###############################################################################
#TSMC Library/IP Product
#Filename: tcb018gbwp7t_6lm.lef
#Technology: CL018G
#Product Type: Standard Cell
#Product Name: tcb018gbwp7t
#Version: 270a
###############################################################################
# 
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
# 
###############################################################################

# DESIGN RULE DOCUMENT: T-018-LO-DR-001 V2.7
#+
#+Note:
#+ 1. Use Capatable to substitute 1DRC defined in LEF header is strongly recommended.
#+
# Resistor & Capacitor are referenced from spice model interconnect table
# The index is "width=minWidth", "Space=Pitch"
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    CAPACITANCE PICOFARADS 10 ;
    CURRENT MILLIAMPS 10000 ;
    VOLTAGE VOLTS 1000 ;
    FREQUENCY MEGAHERTZ 10 ;
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER POLY1
    TYPE MASTERSLICE ;
END POLY1

LAYER POLY2
    TYPE MASTERSLICE ;
END POLY2

LAYER CONT
    TYPE CUT ;
END CONT

LAYER METAL1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    OFFSET	0.280 ;
    PITCH	0.560 ;
    WIDTH	0.230 ;
    SPACING	0.230 ;
    AREA	0.202 ;
    THICKNESS	0.530 ;
    HEIGHT	1.100 ;
    MINIMUMDENSITY	30 ;
    SPACING 0.600 RANGE 10.001 200.0 ;
 
    ANTENNASIDEAREARATIO	400.000000 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.2029 400 ) ( 0.203 2281.2 ) ( 0.5 2400 ) ( 1 2600 ) ( 1.5 2800 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
        WIDTH           0.230   1.000 ;
        TABLEENTRIES    1.000   1.000 ;
    ACCURRENTDENSITY    RMS
    FREQUENCY	500 ;
        WIDTH           0.230   1.000 ;
        TABLEENTRIES    8.000   8.000 ;
    ACCURRENTDENSITY    PEAK
    FREQUENCY	500 ;
        WIDTH           0.230   1.000 ;
        TABLEENTRIES    28.284   28.284 ;
    DCCURRENTDENSITY	AVERAGE
        WIDTH           0.230   1.000 ;
        TABLEENTRIES    1.000   1.000 ;

    RESISTANCE RPERSQ 0.0780000000 ;
    CAPACITANCE CPERSQDIST 0.0000473913 ;
    EDGECAPACITANCE 0.0000640000 ;
END METAL1

LAYER VIA12
    TYPE CUT ;
    SPACING	0.260 ;
 
    ANTENNAAREARATIO	20.000000 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.2029 20 ) ( 0.203 91.916 ) ( 0.5 116.665 ) ( 1 158.33 ) ( 1.5 199.995 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
    TABLEENTRIES	4.14201183 ;
END VIA12

LAYER METAL2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    OFFSET	0.280 ;
    PITCH	0.560 ;
    WIDTH	0.280 ;
    SPACING	0.280 ;
    AREA	0.202 ;
    THICKNESS	0.530 ;
    HEIGHT	2.480 ;
    MINIMUMDENSITY	30 ;
    SPACING 0.600 RANGE 10.001 200.0 ;

    ANTENNASIDEAREARATIO	400.000000 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.2029 400 ) ( 0.203 2281.2 ) ( 0.5 2400 ) ( 1 2600 ) ( 1.5 2800 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;
    ACCURRENTDENSITY    RMS
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    4.000   4.000 ;        
    ACCURRENTDENSITY    PEAK
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    28.284   28.284 ;
    DCCURRENTDENSITY AVERAGE
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;

    RESISTANCE RPERSQ 0.0780000000 ;
    CAPACITANCE CPERSQDIST 0.0000396429 ;
    EDGECAPACITANCE 0.0000683000 ;
END METAL2

LAYER VIA23
    TYPE CUT ;
    SPACING	0.260 ;
 
    ANTENNAAREARATIO	20.000000 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.2029 20 ) ( 0.203 91.916 ) ( 0.5 116.665 ) ( 1 158.33 ) ( 1.5 199.995 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
    TABLEENTRIES	4.14201183 ;
END VIA23

LAYER METAL3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    OFFSET	0.280 ;
    PITCH	0.560 ;
    WIDTH	0.280 ;
    SPACING	0.280 ;
    AREA	0.202 ;
    THICKNESS	0.530 ;
    HEIGHT	3.860 ;
    MINIMUMDENSITY	30 ;
    SPACING 0.600 RANGE 10.001 200.0 ;

    ANTENNASIDEAREARATIO	400.000000 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.2029 400 ) ( 0.203 2281.2 ) ( 0.5 2400 ) ( 1 2600 ) ( 1.5 2800 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;
    ACCURRENTDENSITY    RMS
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    4.000   4.000 ;
    ACCURRENTDENSITY    PEAK
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    28.284   28.284 ;
    DCCURRENTDENSITY AVERAGE
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;

    RESISTANCE RPERSQ 0.0780000000 ;
    CAPACITANCE CPERSQDIST 0.0000396429 ;
    EDGECAPACITANCE 0.0000682000 ;
END METAL3

LAYER VIA34
    TYPE CUT ;
    SPACING	0.260 ;
 
    ANTENNAAREARATIO	20.000000 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.2029 20 ) ( 0.203 91.916 ) ( 0.5 116.665 ) ( 1 158.33 ) ( 1.5 199.995 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
    TABLEENTRIES	4.14201183 ;
END VIA34

LAYER METAL4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    OFFSET	0.280 ;
    PITCH	0.560 ;
    WIDTH	0.280 ;
    SPACING	0.280 ;
    AREA	0.202 ;
    THICKNESS	0.530 ;
    HEIGHT	5.240 ;
    MINIMUMDENSITY	30 ;
    SPACING 0.600 RANGE 10.001 200.0 ;

    ANTENNASIDEAREARATIO	400.000000 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.2029 400 ) ( 0.203 2281.2 ) ( 0.5 2400 ) ( 1 2600 ) ( 1.5 2800 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;
    ACCURRENTDENSITY    RMS
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    4.000   4.000 ;        
    ACCURRENTDENSITY    PEAK
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    28.284   28.284 ;
    DCCURRENTDENSITY AVERAGE
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;

    RESISTANCE RPERSQ 0.0780000000 ;
    CAPACITANCE CPERSQDIST 0.0000396429 ;
    EDGECAPACITANCE 0.0000682000 ;
END METAL4

LAYER VIA45
    TYPE CUT ;
    SPACING	0.260 ;
 
    ANTENNAAREARATIO	20.000000 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.2029 20 ) ( 0.203 91.916 ) ( 0.5 116.665 ) ( 1 158.33 ) ( 1.5 199.995 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
    TABLEENTRIES	4.14201183 ;
END VIA45

LAYER METAL5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    OFFSET	0.280 ;
    PITCH	0.560 ;
    WIDTH	0.280 ;
    SPACING	0.280 ;
    AREA	0.202 ;
    THICKNESS	0.530 ;
    HEIGHT	6.620 ;
    MINIMUMDENSITY	30 ;
    SPACING 0.600 RANGE 10.001 200.0 ;

    ANTENNASIDEAREARATIO	400.000000 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.2029 400 ) ( 0.203 2281.2 ) ( 0.5 2400 ) ( 1 2600 ) ( 1.5 2800 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;
    ACCURRENTDENSITY    RMS
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    4.000   4.000 ;        
    ACCURRENTDENSITY    PEAK
    FREQUENCY	500 ;
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    28.284   28.284 ;
    DCCURRENTDENSITY AVERAGE
        WIDTH           0.280   1.000 ;
        TABLEENTRIES    1.000   1.000 ;

    RESISTANCE RPERSQ 0.0780000000 ;
    CAPACITANCE CPERSQDIST 0.0000396429 ;
    EDGECAPACITANCE 0.0000680000 ;
END METAL5

LAYER VIA56
    TYPE CUT ;
    SPACING	0.350 ;
 
    ANTENNAAREARATIO	20.000000 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.2029 20 ) ( 0.203 91.916 ) ( 0.5 116.665 ) ( 1 158.33 ) ( 1.5 199.995 ) ) ;
    
    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
    TABLEENTRIES	5.44753086 ;
END VIA56

LAYER METAL6
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    OFFSET	0.280 ;
    PITCH	0.900 ;
    WIDTH	0.440 ;
    SPACING	0.460 ;
    AREA	0.562 ;
    THICKNESS	0.990 ;
    HEIGHT	8.150 ;
    MINIMUMDENSITY	30 ;
    SPACING 0.600 RANGE 10.001 200.0 ;

    ANTENNASIDEAREARATIO	400.000000 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.2029 400 ) ( 0.203 31624 ) ( 0.5 34000 ) ( 1 38000 ) ( 1.5 42000 ) ) ;

    ACCURRENTDENSITY    AVERAGE
    FREQUENCY	500 ;
        WIDTH           0.440   1.000 ;
        TABLEENTRIES    1.600   1.600 ;
    ACCURRENTDENSITY    RMS
    FREQUENCY	500 ;
        WIDTH           0.440   1.000 ;
        TABLEENTRIES    8.000   8.000 ;
    ACCURRENTDENSITY    PEAK
    FREQUENCY	500 ;
        WIDTH           0.440   1.000 ;
        TABLEENTRIES    56.568   56.568 ;
    DCCURRENTDENSITY AVERAGE
        WIDTH           0.440   1.000 ;
        TABLEENTRIES    1.600   1.600 ;

    RESISTANCE RPERSQ 0.0360000000 ;
    CAPACITANCE CPERSQDIST 0.0000340909 ;
    EDGECAPACITANCE 0.0000784000 ;
END METAL6

LAYER OVERLAP
    TYPE OVERLAP ;
END OVERLAP

VIA VIA12_HV DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL1 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA12 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL2 ;
        RECT -0.140 -0.190 0.140 0.190 ;
END VIA12_HV

VIA VIA12_VH DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL1 ;
        RECT -0.140 -0.190 0.140 0.190 ;
    LAYER VIA12 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL2 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA12_VH

VIA VIA12_HH DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL1 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA12 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL2 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA12_HH
                   
VIA VIA12_VV DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL1 ;
        RECT -0.140 -0.190 0.140 0.190 ;
    LAYER VIA12 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL2 ;
        RECT -0.140 -0.190 0.140 0.190 ;
END VIA12_VV
                   
VIA VIA2 DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL2 ;
        RECT -0.140 -0.190 0.140 0.190 ;
    LAYER VIA23 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA2

VIA VIA2NORTH DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL2 ;
        RECT -0.140 -0.190 0.140 0.535 ;
    LAYER VIA23 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA2NORTH
                   
VIA VIA2SOUTH DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL2 ;
        RECT -0.140 -0.535 0.140 0.190 ;
    LAYER VIA23 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA2SOUTH

VIA VIA3 DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.190 0.140 ;
    LAYER VIA34 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL4 ;
        RECT -0.140 -0.190 0.140 0.190 ;
END VIA3

VIA VIA3EAST DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL3 ;
        RECT -0.190 -0.140 0.535 0.140 ;
    LAYER VIA34 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL4 ;
        RECT -0.140 -0.190 0.140 0.190 ;
END VIA3EAST
                   
VIA VIA3WEST DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL3 ;
        RECT -0.535 -0.140 0.190 0.140 ;
    LAYER VIA34 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL4 ;
        RECT -0.140 -0.190 0.140 0.190 ;
END VIA3WEST

VIA VIA4 DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL4 ;
        RECT -0.140 -0.190 0.140 0.190 ;
    LAYER VIA45 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL5 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA4

VIA VIA4NORTH DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL4 ;
        RECT -0.140 -0.190 0.140 0.535 ;
    LAYER VIA45 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL5 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA4NORTH
                   
VIA VIA4SOUTH DEFAULT
    RESISTANCE 6.4000000000 ;
    LAYER METAL4 ;
        RECT -0.140 -0.535 0.140 0.190 ;
    LAYER VIA45 ;
        RECT -0.130 -0.130 0.130 0.130 ;
    LAYER METAL5 ;
        RECT -0.190 -0.140 0.190 0.140 ;
END VIA4SOUTH

VIA VIA5 DEFAULT
    RESISTANCE 2.5400000000 ;
    LAYER METAL5 ;
        RECT -0.240 -0.190 0.240 0.190 ;
    LAYER VIA56 ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER METAL6 ;
        RECT -0.270 -0.270 0.270 0.270 ;
END VIA5

VIA VIA5EAST DEFAULT
    RESISTANCE 2.5400000000 ;
    LAYER METAL5 ;
        RECT -0.240 -0.190 0.295 0.190 ;
    LAYER VIA56 ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER METAL6 ;
        RECT -0.270 -0.270 0.270 0.270 ;
END VIA5EAST
                   
VIA VIA5WEST DEFAULT
    RESISTANCE 2.5400000000 ;
    LAYER METAL5 ;
        RECT -0.295 -0.190 0.240 0.190 ;
    LAYER VIA56 ;
        RECT -0.180 -0.180 0.180 0.180 ;
    LAYER METAL6 ;
        RECT -0.270 -0.270 0.270 0.270 ;
END VIA5WEST

VIARULE VIAGEN12 GENERATE
    LAYER METAL1 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER METAL2 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER VIA12 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END VIAGEN12        

VIARULE VIAGEN23 GENERATE
    LAYER METAL2 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER METAL3 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER VIA23 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END VIAGEN23

VIARULE VIAGEN34 GENERATE
    LAYER METAL3 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER METAL4 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER VIA34 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END VIAGEN34

VIARULE VIAGEN45 GENERATE
    LAYER METAL4 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER METAL5 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER VIA45 ;
        RECT -0.130 -0.130 0.130 0.130 ;
        SPACING 0.520 BY 0.520 ;
END VIAGEN45

VIARULE VIAGEN56 GENERATE
    LAYER METAL5 ;
        ENCLOSURE 0.060 0.010 ;
    LAYER METAL6 ;
        ENCLOSURE 0.090 0.090 ;
    LAYER VIA56 ;
        RECT -0.180 -0.180 0.180 0.180 ;
        SPACING 0.710 BY 0.710 ;
END VIAGEN56

SITE core7T
    CLASS CORE ;
    SYMMETRY Y  ;
    SIZE 0.560 BY 3.920 ;
END core7T

SITE bcore7T
    CLASS CORE ;
    SYMMETRY Y  ;
    SIZE 0.560 BY 7.840 ;
END bcore7T

SITE bcoreExt7T
    SIZE 0.560 BY 7.840 ;
    CLASS CORE ;
END bcoreExt7T

SITE ccore7T
    CLASS CORE ;
    SYMMETRY Y  ;
    SIZE 0.560 BY 11.760 ;
END ccore7T

SITE dcore7T
    CLASS CORE ;
    SYMMETRY Y  ;
    SIZE 0.560 BY 15.680 ;
END dcore7T

SITE gacore7T
    CLASS CORE ;
    SYMMETRY Y  ;
    SIZE 2.240 BY 3.920 ;
END gacore7T

MACRO AN2D0BWP7T
    CLASS CORE ;
    FOREIGN AN2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 0.580 2.660 2.715 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        RECT  1.145 1.480 1.260 1.820 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.420 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 -0.235 2.800 0.235 ;
        RECT  1.540 -0.235 1.920 0.870 ;
        RECT  0.000 -0.235 1.540 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.815 3.685 2.800 4.155 ;
        RECT  1.390 3.405 1.815 4.155 ;
        RECT  0.520 3.685 1.390 4.155 ;
        RECT  0.170 3.400 0.520 4.155 ;
        RECT  0.000 3.685 0.170 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.840 1.480 2.100 2.695 ;
        RECT  0.915 2.455 1.840 2.695 ;
        RECT  0.685 0.630 0.915 2.695 ;
        RECT  0.180 0.630 0.685 0.870 ;
    END
END AN2D0BWP7T

MACRO AN2D1BWP7T
    CLASS CORE ;
    FOREIGN AN2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 0.465 2.660 3.300 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.655 0.455 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 -0.235 2.800 0.235 ;
        RECT  1.485 -0.235 1.825 0.720 ;
        RECT  0.000 -0.235 1.485 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 3.685 2.800 4.155 ;
        RECT  1.560 3.015 1.900 4.155 ;
        RECT  0.525 3.685 1.560 4.155 ;
        RECT  0.185 3.450 0.525 4.155 ;
        RECT  0.000 3.685 0.185 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.855 1.605 2.085 2.680 ;
        RECT  0.945 2.450 1.855 2.680 ;
        RECT  0.685 0.470 0.945 2.680 ;
        RECT  0.180 0.470 0.685 0.700 ;
    END
END AN2D1BWP7T

MACRO AN2D2BWP7T
    CLASS CORE ;
    FOREIGN AN2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.475 ;
        RECT  2.745 1.210 2.940 1.655 ;
        RECT  2.745 2.245 2.940 2.475 ;
        RECT  2.515 0.475 2.745 1.655 ;
        RECT  2.515 2.245 2.745 3.375 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 1.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.630 0.460 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 -0.235 3.920 0.235 ;
        RECT  3.160 -0.235 3.540 0.890 ;
        RECT  2.110 -0.235 3.160 0.235 ;
        RECT  1.730 -0.235 2.110 0.800 ;
        RECT  0.000 -0.235 1.730 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 3.685 3.920 4.155 ;
        RECT  3.160 2.725 3.540 4.155 ;
        RECT  2.115 3.685 3.160 4.155 ;
        RECT  1.730 2.900 2.115 4.155 ;
        RECT  0.670 3.685 1.730 4.155 ;
        RECT  0.290 3.025 0.670 4.155 ;
        RECT  0.000 3.685 0.290 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.010 1.075 2.250 2.670 ;
        RECT  0.585 1.075 2.010 1.305 ;
        RECT  1.305 2.430 2.010 2.670 ;
        RECT  1.075 2.430 1.305 3.350 ;
        RECT  0.355 0.465 0.585 1.305 ;
    END
END AN2D2BWP7T

MACRO AN2D4BWP7T
    CLASS CORE ;
    FOREIGN AN2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.535 0.495 5.770 3.335 ;
        RECT  4.870 1.050 5.535 2.605 ;
        RECT  4.265 1.050 4.870 1.340 ;
        RECT  4.265 2.255 4.870 2.605 ;
        RECT  4.035 0.485 4.265 1.340 ;
        RECT  4.035 2.255 4.265 3.335 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.785 1.660 3.015 2.370 ;
        RECT  0.980 2.140 2.785 2.370 ;
        RECT  0.700 1.705 0.980 2.370 ;
        RECT  0.140 1.705 0.700 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.635 2.360 1.865 ;
        RECT  1.260 0.650 1.540 1.865 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.495 -0.235 6.720 0.235 ;
        RECT  6.250 -0.235 6.495 1.300 ;
        RECT  5.100 -0.235 6.250 0.235 ;
        RECT  4.720 -0.235 5.100 0.785 ;
        RECT  3.600 -0.235 4.720 0.235 ;
        RECT  3.240 -0.235 3.600 0.785 ;
        RECT  0.470 -0.235 3.240 0.235 ;
        RECT  0.230 -0.235 0.470 1.240 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.510 3.685 6.720 4.155 ;
        RECT  6.225 2.255 6.510 4.155 ;
        RECT  5.090 3.685 6.225 4.155 ;
        RECT  4.710 3.015 5.090 4.155 ;
        RECT  3.595 3.685 4.710 4.155 ;
        RECT  3.215 3.155 3.595 4.155 ;
        RECT  2.110 3.685 3.215 4.155 ;
        RECT  1.730 3.155 2.110 4.155 ;
        RECT  0.480 3.685 1.730 4.155 ;
        RECT  0.220 2.460 0.480 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.265 1.050 4.670 1.340 ;
        RECT  4.265 2.255 4.670 2.605 ;
        RECT  4.035 0.485 4.265 1.340 ;
        RECT  4.035 2.255 4.265 3.335 ;
        RECT  3.635 1.660 4.550 1.920 ;
        RECT  3.405 1.090 3.635 2.900 ;
        RECT  2.015 1.090 3.405 1.320 ;
        RECT  2.785 2.610 3.405 2.900 ;
        RECT  2.555 2.610 2.785 3.450 ;
        RECT  1.245 2.610 2.555 2.900 ;
        RECT  1.785 0.495 2.015 1.320 ;
        RECT  1.015 2.610 1.245 3.450 ;
    END
END AN2D4BWP7T

MACRO AN2XD1BWP7T
    CLASS CORE ;
    FOREIGN AN2XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1968 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.020 3.225 2.480 ;
        RECT  2.930 1.020 2.940 1.305 ;
        RECT  2.930 2.245 2.940 2.480 ;
        RECT  2.700 0.495 2.930 1.305 ;
        RECT  2.700 2.245 2.930 3.365 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.610 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.670 0.455 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.155 -0.235 3.360 0.235 ;
        RECT  1.905 -0.235 2.155 1.270 ;
        RECT  0.000 -0.235 1.905 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.225 3.685 3.360 4.155 ;
        RECT  1.845 2.990 2.225 4.155 ;
        RECT  0.595 3.685 1.845 4.155 ;
        RECT  0.215 3.050 0.595 4.155 ;
        RECT  0.000 3.685 0.215 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.220 1.655 2.450 2.740 ;
        RECT  1.300 2.465 2.220 2.740 ;
        RECT  1.070 2.465 1.300 3.230 ;
        RECT  1.015 2.465 1.070 2.740 ;
        RECT  0.785 1.130 1.015 2.740 ;
        RECT  0.530 1.130 0.785 1.360 ;
        RECT  0.285 0.485 0.530 1.360 ;
    END
END AN2XD1BWP7T

MACRO AN3D0BWP7T
    CLASS CORE ;
    FOREIGN AN3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 0.570 3.220 2.710 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.160 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 0.650 1.540 1.590 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.460 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.530 -0.235 3.360 0.235 ;
        RECT  2.070 -0.235 2.530 0.870 ;
        RECT  0.000 -0.235 2.070 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.195 3.685 3.360 4.155 ;
        RECT  1.835 3.415 2.195 4.155 ;
        RECT  1.100 3.685 1.835 4.155 ;
        RECT  0.720 3.415 1.100 4.155 ;
        RECT  0.000 3.685 0.720 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.665 3.135 2.980 3.365 ;
        RECT  2.435 2.435 2.665 3.365 ;
        RECT  0.930 2.435 2.435 2.675 ;
        RECT  0.700 0.635 0.930 2.675 ;
        RECT  0.180 0.635 0.700 0.875 ;
        RECT  0.180 2.435 0.700 2.675 ;
    END
END AN3D0BWP7T

MACRO AN3D1BWP7T
    CLASS CORE ;
    FOREIGN AN3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.485 3.220 3.425 ;
        RECT  2.895 0.485 2.940 1.305 ;
        RECT  2.895 2.375 2.940 3.425 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 1.210 2.100 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.170 0.650 1.540 1.590 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.475 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.445 -0.235 3.360 0.235 ;
        RECT  2.065 -0.235 2.445 0.750 ;
        RECT  0.000 -0.235 2.065 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.410 3.685 3.360 4.155 ;
        RECT  2.065 3.410 2.410 4.155 ;
        RECT  1.135 3.685 2.065 4.155 ;
        RECT  0.720 3.415 1.135 4.155 ;
        RECT  0.000 3.685 0.720 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.610 1.605 2.710 1.945 ;
        RECT  2.350 1.605 2.610 2.720 ;
        RECT  0.935 2.480 2.350 2.720 ;
        RECT  0.705 0.470 0.935 2.720 ;
        RECT  0.180 0.470 0.705 0.720 ;
        RECT  0.180 2.480 0.705 2.720 ;
    END
END AN3D1BWP7T

MACRO AN3D2BWP7T
    CLASS CORE ;
    FOREIGN AN3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.100 3.780 2.455 ;
        RECT  3.385 1.100 3.500 1.330 ;
        RECT  3.385 2.225 3.500 2.455 ;
        RECT  3.155 0.475 3.385 1.330 ;
        RECT  3.155 2.225 3.385 3.405 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.660 2.185 2.150 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 0.650 1.560 1.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.460 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 -0.235 4.480 0.235 ;
        RECT  4.015 -0.235 4.245 1.265 ;
        RECT  2.740 -0.235 4.015 0.235 ;
        RECT  2.360 -0.235 2.740 1.195 ;
        RECT  0.000 -0.235 2.360 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 3.685 4.480 4.155 ;
        RECT  4.015 2.245 4.245 4.155 ;
        RECT  2.745 3.685 4.015 4.155 ;
        RECT  2.365 3.155 2.745 4.155 ;
        RECT  1.300 3.685 2.365 4.155 ;
        RECT  0.920 3.155 1.300 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.890 1.660 3.200 1.890 ;
        RECT  2.660 1.660 2.890 2.780 ;
        RECT  1.945 2.550 2.660 2.780 ;
        RECT  1.715 2.550 1.945 3.305 ;
        RECT  0.970 2.550 1.715 2.780 ;
        RECT  0.730 0.665 0.970 2.780 ;
        RECT  0.210 0.665 0.730 0.895 ;
        RECT  0.505 2.550 0.730 2.780 ;
        RECT  0.275 2.550 0.505 3.360 ;
    END
END AN3D2BWP7T

MACRO AN3D4BWP7T
    CLASS CORE ;
    FOREIGN AN3D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.090 0.495 7.375 1.460 ;
        RECT  7.090 2.255 7.375 3.430 ;
        RECT  6.890 1.060 7.090 1.460 ;
        RECT  6.890 2.255 7.090 2.605 ;
        RECT  5.990 1.060 6.890 2.605 ;
        RECT  5.790 1.060 5.990 1.410 ;
        RECT  5.790 2.255 5.990 2.605 ;
        RECT  5.520 0.495 5.790 1.410 ;
        RECT  5.520 2.255 5.790 3.430 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.280 1.190 4.510 1.980 ;
        RECT  0.465 1.190 4.280 1.420 ;
        RECT  0.140 1.190 0.465 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 1.680 3.750 2.710 ;
        RECT  1.540 2.475 3.520 2.710 ;
        RECT  1.260 1.735 1.540 2.710 ;
        RECT  1.145 1.735 1.260 1.980 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.730 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.070 -0.235 8.400 0.235 ;
        RECT  7.840 -0.235 8.070 1.290 ;
        RECT  6.660 -0.235 7.840 0.235 ;
        RECT  6.280 -0.235 6.660 0.790 ;
        RECT  4.995 -0.235 6.280 0.235 ;
        RECT  4.590 -0.235 4.995 0.470 ;
        RECT  0.540 -0.235 4.590 0.235 ;
        RECT  0.160 -0.235 0.540 0.870 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.070 3.685 8.400 4.155 ;
        RECT  7.840 2.245 8.070 4.155 ;
        RECT  6.650 3.685 7.840 4.155 ;
        RECT  6.270 3.090 6.650 4.155 ;
        RECT  5.085 3.685 6.270 4.155 ;
        RECT  4.705 2.940 5.085 4.155 ;
        RECT  3.545 3.685 4.705 4.155 ;
        RECT  3.185 3.450 3.545 4.155 ;
        RECT  2.045 3.685 3.185 4.155 ;
        RECT  1.655 3.440 2.045 4.155 ;
        RECT  0.465 3.685 1.655 4.155 ;
        RECT  0.235 2.405 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.090 0.495 7.375 1.460 ;
        RECT  7.090 2.255 7.375 3.430 ;
        RECT  5.520 0.495 5.790 1.410 ;
        RECT  5.520 2.255 5.790 3.430 ;
        RECT  4.985 1.735 5.685 1.965 ;
        RECT  4.755 0.700 4.985 2.660 ;
        RECT  2.405 0.700 4.755 0.955 ;
        RECT  4.355 2.430 4.755 2.660 ;
        RECT  4.125 2.430 4.355 3.195 ;
        RECT  0.885 2.940 4.125 3.195 ;
    END
END AN3D4BWP7T

MACRO AN3XD1BWP7T
    CLASS CORE ;
    FOREIGN AN3XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.4220 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.940 3.780 2.670 ;
        RECT  3.450 0.940 3.500 1.305 ;
        RECT  3.450 2.250 3.500 2.670 ;
        RECT  3.220 0.485 3.450 1.305 ;
        RECT  3.220 2.250 3.450 3.360 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.175 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 0.650 1.540 2.020 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.520 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.665 -0.235 3.920 0.235 ;
        RECT  2.285 -0.235 2.665 0.940 ;
        RECT  0.000 -0.235 2.285 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 3.685 3.920 4.155 ;
        RECT  2.365 3.155 2.745 4.155 ;
        RECT  1.290 3.685 2.365 4.155 ;
        RECT  0.910 3.155 1.290 4.155 ;
        RECT  0.000 3.685 0.910 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.680 1.660 2.910 2.695 ;
        RECT  1.940 2.465 2.680 2.695 ;
        RECT  1.710 2.465 1.940 3.395 ;
        RECT  0.990 2.465 1.710 2.695 ;
        RECT  0.760 0.685 0.990 2.695 ;
        RECT  0.215 0.685 0.760 0.915 ;
        RECT  0.500 2.465 0.760 2.695 ;
        RECT  0.270 2.465 0.500 3.395 ;
    END
END AN3XD1BWP7T

MACRO AN4D0BWP7T
    CLASS CORE ;
    FOREIGN AN4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5797 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.465 3.780 2.735 ;
        RECT  3.455 0.465 3.500 0.820 ;
        RECT  3.455 2.310 3.500 2.735 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 1.210 2.660 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 1.055 2.100 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        RECT  1.140 1.680 1.260 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 -0.235 3.920 0.235 ;
        RECT  2.605 -0.235 3.065 0.715 ;
        RECT  0.000 -0.235 2.605 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 3.685 3.920 4.155 ;
        RECT  2.580 3.400 2.820 4.155 ;
        RECT  2.350 3.685 2.580 4.155 ;
        RECT  2.110 3.400 2.350 4.155 ;
        RECT  1.880 3.685 2.110 4.155 ;
        RECT  1.640 3.400 1.880 4.155 ;
        RECT  1.410 3.685 1.640 4.155 ;
        RECT  1.170 3.400 1.410 4.155 ;
        RECT  0.940 3.685 1.170 4.155 ;
        RECT  0.700 3.400 0.940 4.155 ;
        RECT  0.470 3.685 0.700 4.155 ;
        RECT  0.230 3.400 0.470 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.190 1.360 3.270 1.705 ;
        RECT  2.960 1.360 3.190 2.705 ;
        RECT  0.910 2.475 2.960 2.705 ;
        RECT  0.680 0.490 0.910 2.705 ;
        RECT  0.180 0.490 0.680 0.720 ;
    END
END AN4D0BWP7T

MACRO AN4D1BWP7T
    CLASS CORE ;
    FOREIGN AN4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1595 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.485 3.780 3.335 ;
        RECT  3.455 0.485 3.500 1.315 ;
        RECT  3.455 2.310 3.500 3.335 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 1.210 2.660 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 1.055 2.100 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        RECT  1.140 1.680 1.260 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 -0.235 3.920 0.235 ;
        RECT  2.605 -0.235 3.065 0.715 ;
        RECT  0.000 -0.235 2.605 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 3.685 3.920 4.155 ;
        RECT  2.580 3.400 2.820 4.155 ;
        RECT  2.350 3.685 2.580 4.155 ;
        RECT  2.110 3.400 2.350 4.155 ;
        RECT  1.880 3.685 2.110 4.155 ;
        RECT  1.640 3.400 1.880 4.155 ;
        RECT  1.410 3.685 1.640 4.155 ;
        RECT  1.170 3.400 1.410 4.155 ;
        RECT  0.940 3.685 1.170 4.155 ;
        RECT  0.700 3.400 0.940 4.155 ;
        RECT  0.470 3.685 0.700 4.155 ;
        RECT  0.230 3.400 0.470 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.190 1.660 3.270 2.005 ;
        RECT  2.960 1.660 3.190 2.705 ;
        RECT  0.910 2.475 2.960 2.705 ;
        RECT  0.680 0.490 0.910 2.705 ;
        RECT  0.180 0.490 0.680 0.720 ;
    END
END AN4D1BWP7T

MACRO AN4D2BWP7T
    CLASS CORE ;
    FOREIGN AN4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 1.170 4.340 2.750 ;
        RECT  4.060 0.495 4.085 3.340 ;
        RECT  3.855 0.495 4.060 1.410 ;
        RECT  3.855 2.480 4.060 3.340 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.700 1.620 2.905 2.190 ;
        RECT  2.380 1.210 2.700 2.190 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.650 2.115 1.915 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 1.210 1.575 2.190 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.630 0.480 2.715 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 -0.235 5.040 0.235 ;
        RECT  4.575 -0.235 4.805 1.300 ;
        RECT  3.445 -0.235 4.575 0.235 ;
        RECT  3.065 -0.235 3.445 1.185 ;
        RECT  0.000 -0.235 3.065 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 3.685 5.040 4.155 ;
        RECT  4.575 2.255 4.805 4.155 ;
        RECT  3.435 3.685 4.575 4.155 ;
        RECT  3.055 3.115 3.435 4.155 ;
        RECT  2.000 3.685 3.055 4.155 ;
        RECT  1.620 3.115 2.000 4.155 ;
        RECT  0.555 3.685 1.620 4.155 ;
        RECT  0.175 3.115 0.555 4.155 ;
        RECT  0.000 3.685 0.175 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.610 1.715 3.780 1.945 ;
        RECT  3.380 1.715 3.610 2.790 ;
        RECT  2.645 2.560 3.380 2.790 ;
        RECT  2.415 2.560 2.645 3.395 ;
        RECT  1.205 2.560 2.415 2.790 ;
        RECT  0.975 2.560 1.205 3.400 ;
        RECT  0.955 2.560 0.975 2.790 ;
        RECT  0.725 1.090 0.955 2.790 ;
        RECT  0.480 1.090 0.725 1.325 ;
        RECT  0.250 0.495 0.480 1.325 ;
    END
END AN4D2BWP7T

MACRO AN4D4BWP7T
    CLASS CORE ;
    FOREIGN AN4D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 0.495 9.130 3.345 ;
        RECT  8.230 0.935 8.895 2.580 ;
        RECT  7.400 0.935 8.230 1.285 ;
        RECT  7.690 2.230 8.230 2.580 ;
        RECT  7.450 2.230 7.690 3.345 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.530 0.860 6.760 1.885 ;
        RECT  6.465 0.860 6.530 1.090 ;
        RECT  6.235 0.465 6.465 1.090 ;
        RECT  0.980 0.465 6.235 0.695 ;
        RECT  0.700 0.465 0.980 2.150 ;
        RECT  0.690 1.475 0.700 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.545 1.780 5.820 2.010 ;
        RECT  5.315 1.385 5.545 2.010 ;
        RECT  3.590 1.385 5.315 1.615 ;
        RECT  3.360 0.925 3.590 1.615 ;
        RECT  1.540 0.925 3.360 1.155 ;
        RECT  1.540 1.485 1.590 1.825 ;
        RECT  1.260 0.925 1.540 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.8298 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.960 1.845 5.085 2.075 ;
        RECT  4.730 1.845 4.960 2.660 ;
        RECT  4.010 2.380 4.730 2.660 ;
        RECT  2.670 2.380 4.010 2.610 ;
        RECT  2.440 1.845 2.670 2.610 ;
        RECT  2.330 1.845 2.440 2.075 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8298 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 1.845 4.300 2.075 ;
        RECT  2.900 1.385 3.130 2.075 ;
        RECT  2.100 1.385 2.900 1.615 ;
        RECT  1.820 1.385 2.100 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.910 -0.235 10.080 0.235 ;
        RECT  9.530 -0.235 9.910 1.215 ;
        RECT  8.485 -0.235 9.530 0.235 ;
        RECT  8.105 -0.235 8.485 0.700 ;
        RECT  6.925 -0.235 8.105 0.235 ;
        RECT  6.695 -0.235 6.925 0.520 ;
        RECT  0.470 -0.235 6.695 0.235 ;
        RECT  0.240 -0.235 0.470 1.240 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.910 3.685 10.080 4.155 ;
        RECT  9.530 2.300 9.910 4.155 ;
        RECT  8.475 3.685 9.530 4.155 ;
        RECT  8.095 3.035 8.475 4.155 ;
        RECT  7.035 3.685 8.095 4.155 ;
        RECT  6.655 3.240 7.035 4.155 ;
        RECT  5.540 3.685 6.655 4.155 ;
        RECT  5.200 3.455 5.540 4.155 ;
        RECT  4.020 3.685 5.200 4.155 ;
        RECT  3.680 3.455 4.020 4.155 ;
        RECT  2.305 3.685 3.680 4.155 ;
        RECT  1.965 3.455 2.305 4.155 ;
        RECT  0.730 3.685 1.965 4.155 ;
        RECT  0.390 2.635 0.730 4.155 ;
        RECT  0.000 3.685 0.390 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.400 0.935 8.030 1.285 ;
        RECT  7.690 2.230 8.030 2.580 ;
        RECT  7.450 2.230 7.690 3.345 ;
        RECT  7.220 1.590 7.540 1.820 ;
        RECT  6.990 1.590 7.220 2.355 ;
        RECT  6.300 2.115 6.990 2.355 ;
        RECT  1.120 2.995 6.060 3.225 ;
        RECT  5.775 0.925 6.005 1.550 ;
        RECT  3.820 0.925 5.775 1.155 ;
        RECT  6.060 1.320 6.300 3.225 ;
        RECT  6.005 1.320 6.060 1.550 ;
    END
END AN4D4BWP7T

MACRO AN4XD1BWP7T
    CLASS CORE ;
    FOREIGN AN4XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.495 4.340 3.365 ;
        RECT  3.955 0.495 4.060 1.305 ;
        RECT  3.955 2.385 4.060 3.365 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.150 ;
        RECT  2.795 1.600 2.940 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.650 2.200 2.040 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.620 0.465 2.750 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 -0.235 4.480 0.235 ;
        RECT  3.115 -0.235 3.495 0.945 ;
        RECT  0.000 -0.235 3.115 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 3.685 4.480 4.155 ;
        RECT  3.140 3.010 3.520 4.155 ;
        RECT  2.040 3.685 3.140 4.155 ;
        RECT  1.660 3.015 2.040 4.155 ;
        RECT  0.580 3.685 1.660 4.155 ;
        RECT  0.200 3.155 0.580 4.155 ;
        RECT  0.000 3.685 0.200 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.475 1.540 3.705 2.750 ;
        RECT  2.705 2.520 3.475 2.750 ;
        RECT  2.475 2.520 2.705 3.360 ;
        RECT  1.245 2.520 2.475 2.750 ;
        RECT  1.015 2.520 1.245 3.360 ;
        RECT  1.000 2.520 1.015 2.750 ;
        RECT  0.770 1.115 1.000 2.750 ;
        RECT  0.505 1.115 0.770 1.345 ;
        RECT  0.275 0.485 0.505 1.345 ;
    END
END AN4XD1BWP7T

MACRO ANTENNABWP7T
    CLASS CORE ;
    FOREIGN ANTENNABWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN I
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 0.620 0.465 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 1.120 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 1.120 4.155 ;
        END
    END VDD
END ANTENNABWP7T

MACRO AO211D0BWP7T
    CLASS CORE ;
    FOREIGN AO211D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 0.735 3.780 3.320 ;
        RECT  3.390 0.735 3.550 0.965 ;
        RECT  3.455 2.330 3.550 3.320 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 2.330 3.220 2.710 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.790 2.710 2.100 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        RECT  1.145 1.795 1.260 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 -0.235 3.920 0.235 ;
        RECT  2.630 -0.235 2.970 0.465 ;
        RECT  1.710 -0.235 2.630 0.235 ;
        RECT  1.370 -0.235 1.710 0.465 ;
        RECT  0.000 -0.235 1.370 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 3.685 3.920 4.155 ;
        RECT  2.680 3.040 3.020 4.155 ;
        RECT  0.000 3.685 2.680 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.090 1.250 3.320 1.960 ;
        RECT  2.345 1.250 3.090 1.480 ;
        RECT  2.115 0.695 2.345 1.480 ;
        RECT  0.910 0.695 2.115 0.925 ;
        RECT  0.910 2.625 1.190 2.855 ;
        RECT  0.680 0.695 0.910 2.855 ;
        RECT  0.180 1.015 0.680 1.245 ;
    END
END AO211D0BWP7T

MACRO AO211D1BWP7T
    CLASS CORE ;
    FOREIGN AO211D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.3391 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 1.070 4.340 2.745 ;
        RECT  4.060 0.495 4.245 3.390 ;
        RECT  4.015 0.495 4.060 1.305 ;
        RECT  4.015 2.330 4.060 3.390 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 1.660 3.240 2.710 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.175 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 1.210 1.590 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.715 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 -0.235 4.480 0.235 ;
        RECT  3.145 -0.235 3.525 0.865 ;
        RECT  1.885 -0.235 3.145 0.235 ;
        RECT  1.535 -0.235 1.885 0.890 ;
        RECT  0.000 -0.235 1.535 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 3.685 4.480 4.155 ;
        RECT  3.115 3.075 3.495 4.155 ;
        RECT  0.000 3.685 3.115 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.700 1.660 3.830 2.000 ;
        RECT  3.470 1.120 3.700 2.000 ;
        RECT  2.665 1.120 3.470 1.360 ;
        RECT  2.435 0.495 2.665 2.735 ;
        RECT  0.930 2.505 2.435 2.735 ;
        RECT  0.220 2.965 2.000 3.195 ;
        RECT  0.700 1.075 0.930 2.735 ;
        RECT  0.505 1.075 0.700 1.305 ;
        RECT  0.275 0.495 0.505 1.305 ;
    END
END AO211D1BWP7T

MACRO AO211D2BWP7T
    CLASS CORE ;
    FOREIGN AO211D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.655 4.340 2.645 ;
        RECT  3.740 0.655 4.060 0.885 ;
        RECT  4.025 2.345 4.060 2.645 ;
        RECT  3.795 2.345 4.025 3.415 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.660 3.220 2.710 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.660 2.170 2.150 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 -0.235 5.040 0.235 ;
        RECT  4.575 -0.235 4.805 1.270 ;
        RECT  3.385 -0.235 4.575 0.235 ;
        RECT  3.005 -0.235 3.385 0.865 ;
        RECT  1.930 -0.235 3.005 0.235 ;
        RECT  1.550 -0.235 1.930 0.915 ;
        RECT  0.000 -0.235 1.550 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 3.685 5.040 4.155 ;
        RECT  4.575 2.245 4.805 4.155 ;
        RECT  3.360 3.685 4.575 4.155 ;
        RECT  2.980 3.025 3.360 4.155 ;
        RECT  0.000 3.685 2.980 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.555 1.120 3.785 2.000 ;
        RECT  2.630 1.120 3.555 1.360 ;
        RECT  2.585 1.120 2.630 2.735 ;
        RECT  2.400 0.495 2.585 2.735 ;
        RECT  2.355 0.495 2.400 1.400 ;
        RECT  0.930 2.505 2.400 2.735 ;
        RECT  0.220 3.025 2.000 3.255 ;
        RECT  0.700 1.050 0.930 2.735 ;
        RECT  0.505 1.050 0.700 1.280 ;
        RECT  0.275 0.470 0.505 1.280 ;
    END
END AO211D2BWP7T

MACRO AO21D0BWP7T
    CLASS CORE ;
    FOREIGN AO21D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.555 3.220 3.000 ;
        RECT  2.840 0.555 2.940 0.785 ;
        RECT  2.840 2.770 2.940 3.000 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.200 2.100 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.460 -0.235 3.360 0.235 ;
        RECT  2.120 -0.235 2.460 0.805 ;
        RECT  0.470 -0.235 2.120 0.235 ;
        RECT  0.230 -0.235 0.470 0.860 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 3.685 3.360 4.155 ;
        RECT  2.105 2.915 2.485 4.155 ;
        RECT  0.000 3.685 2.105 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.415 1.950 2.645 2.610 ;
        RECT  1.055 2.380 2.415 2.610 ;
        RECT  0.975 0.615 1.740 0.845 ;
        RECT  0.975 2.380 1.055 3.040 ;
        RECT  0.825 0.615 0.975 3.040 ;
        RECT  0.745 0.615 0.825 2.610 ;
    END
END AO21D0BWP7T

MACRO AO21D1BWP7T
    CLASS CORE ;
    FOREIGN AO21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 1.210 3.780 2.710 ;
        RECT  3.500 0.495 3.625 3.385 ;
        RECT  3.395 0.495 3.500 1.510 ;
        RECT  3.395 2.345 3.500 3.385 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.660 2.305 2.150 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.590 0.515 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 -0.235 3.920 0.235 ;
        RECT  2.545 -0.235 2.925 1.190 ;
        RECT  0.545 -0.235 2.545 0.235 ;
        RECT  0.165 -0.235 0.545 1.245 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 3.685 3.920 4.155 ;
        RECT  2.545 3.005 2.925 4.155 ;
        RECT  0.000 3.685 2.545 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.875 1.660 3.105 2.705 ;
        RECT  1.005 2.475 2.875 2.705 ;
        RECT  1.005 0.665 2.065 0.895 ;
        RECT  0.220 3.045 2.065 3.275 ;
        RECT  0.775 0.665 1.005 2.705 ;
    END
END AO21D1BWP7T

MACRO AO21D2BWP7T
    CLASS CORE ;
    FOREIGN AO21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.170 3.780 2.610 ;
        RECT  3.465 1.170 3.500 1.400 ;
        RECT  3.465 2.380 3.500 2.610 ;
        RECT  3.235 0.465 3.465 1.400 ;
        RECT  3.235 2.380 3.465 3.435 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.660 2.175 2.710 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 -0.235 4.480 0.235 ;
        RECT  4.015 -0.235 4.245 1.245 ;
        RECT  2.730 -0.235 4.015 0.235 ;
        RECT  2.350 -0.235 2.730 0.845 ;
        RECT  0.550 -0.235 2.350 0.235 ;
        RECT  0.170 -0.235 0.550 0.885 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 3.685 4.480 4.155 ;
        RECT  4.015 2.250 4.245 4.155 ;
        RECT  2.785 3.685 4.015 4.155 ;
        RECT  2.405 2.305 2.785 4.155 ;
        RECT  0.000 3.685 2.405 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.675 1.100 2.905 2.000 ;
        RECT  2.120 1.100 2.675 1.330 ;
        RECT  1.890 0.590 2.120 1.330 ;
        RECT  0.505 3.145 2.010 3.375 ;
        RECT  1.010 0.590 1.890 0.820 ;
        RECT  1.010 2.635 1.280 2.865 ;
        RECT  0.780 0.590 1.010 2.865 ;
        RECT  0.275 2.490 0.505 3.375 ;
    END
END AO21D2BWP7T

MACRO AO221D0BWP7T
    CLASS CORE ;
    FOREIGN AO221D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 0.615 4.900 3.045 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.465 0.470 1.805 ;
        RECT  0.140 0.650 0.420 1.805 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.210 3.220 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.220 1.770 2.660 2.150 ;
        RECT  1.820 1.585 2.220 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.540 2.245 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 -0.235 5.040 0.235 ;
        RECT  3.735 -0.235 4.110 0.465 ;
        RECT  2.200 -0.235 3.735 0.235 ;
        RECT  1.820 -0.235 2.200 0.845 ;
        RECT  0.000 -0.235 1.820 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.165 3.685 5.040 4.155 ;
        RECT  3.785 2.915 4.165 4.155 ;
        RECT  0.000 3.685 3.785 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.095 0.695 4.325 2.685 ;
        RECT  2.660 0.695 4.095 0.925 ;
        RECT  1.980 2.455 4.095 2.685 ;
        RECT  3.080 2.915 3.420 3.340 ;
        RECT  0.485 3.110 3.080 3.340 ;
        RECT  2.430 0.695 2.660 1.305 ;
        RECT  0.920 1.075 2.430 1.305 ;
        RECT  1.635 2.455 1.980 2.880 ;
        RECT  0.690 0.830 0.920 1.305 ;
        RECT  0.255 2.720 0.485 3.340 ;
    END
END AO221D0BWP7T

MACRO AO221D1BWP7T
    CLASS CORE ;
    FOREIGN AO221D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 0.495 5.460 3.430 ;
        RECT  5.135 0.495 5.180 1.325 ;
        RECT  5.130 2.405 5.180 3.430 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.050 1.680 4.340 2.710 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.260 2.770 2.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.680 3.780 2.710 ;
        RECT  3.375 1.680 3.500 2.020 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.745 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.730 -0.235 5.600 0.235 ;
        RECT  4.350 -0.235 4.730 0.675 ;
        RECT  2.565 -0.235 4.350 0.235 ;
        RECT  2.190 -0.235 2.565 0.560 ;
        RECT  0.550 -0.235 2.190 0.235 ;
        RECT  0.170 -0.235 0.550 0.930 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.730 3.685 5.600 4.155 ;
        RECT  4.330 3.025 4.730 4.155 ;
        RECT  0.000 3.685 4.330 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.885 1.660 4.950 2.000 ;
        RECT  4.655 1.075 4.885 2.000 ;
        RECT  3.880 1.075 4.655 1.305 ;
        RECT  2.195 3.155 3.980 3.385 ;
        RECT  3.650 0.495 3.880 1.305 ;
        RECT  1.825 0.800 3.650 1.030 ;
        RECT  1.905 2.405 3.260 2.635 ;
        RECT  1.675 2.405 1.905 3.385 ;
        RECT  1.595 0.800 1.825 1.215 ;
        RECT  0.465 3.155 1.675 3.385 ;
        RECT  1.005 0.985 1.595 1.215 ;
        RECT  1.005 2.575 1.240 2.805 ;
        RECT  0.775 0.985 1.005 2.805 ;
        RECT  0.235 2.490 0.465 3.385 ;
    END
END AO221D1BWP7T

MACRO AO221D2BWP7T
    CLASS CORE ;
    FOREIGN AO221D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.765 1.210 6.020 2.600 ;
        RECT  5.740 0.495 5.765 3.365 ;
        RECT  5.535 0.495 5.740 1.440 ;
        RECT  5.535 2.370 5.740 3.365 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.660 4.675 2.000 ;
        RECT  4.060 1.660 4.340 2.710 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.745 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.485 1.210 3.780 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.460 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.730 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 -0.235 6.720 0.235 ;
        RECT  6.255 -0.235 6.485 1.200 ;
        RECT  5.120 -0.235 6.255 0.235 ;
        RECT  4.740 -0.235 5.120 0.785 ;
        RECT  2.735 -0.235 4.740 0.235 ;
        RECT  2.355 -0.235 2.735 0.785 ;
        RECT  0.575 -0.235 2.355 0.235 ;
        RECT  0.195 -0.235 0.575 0.825 ;
        RECT  0.000 -0.235 0.195 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 3.685 6.720 4.155 ;
        RECT  6.255 2.255 6.485 4.155 ;
        RECT  4.985 3.685 6.255 4.155 ;
        RECT  4.755 2.250 4.985 4.155 ;
        RECT  0.000 3.685 4.755 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.245 1.735 5.500 1.965 ;
        RECT  5.015 1.045 5.245 1.965 ;
        RECT  4.370 1.045 5.015 1.275 ;
        RECT  4.130 0.685 4.370 1.275 ;
        RECT  2.470 3.065 4.265 3.295 ;
        RECT  3.250 0.685 4.130 0.915 ;
        RECT  1.945 2.435 3.555 2.665 ;
        RECT  3.020 0.685 3.250 1.250 ;
        RECT  1.825 1.020 3.020 1.250 ;
        RECT  1.715 2.435 1.945 3.430 ;
        RECT  1.595 0.490 1.825 1.250 ;
        RECT  0.505 3.190 1.715 3.430 ;
        RECT  0.970 1.015 1.595 1.250 ;
        RECT  0.970 2.670 1.280 2.900 ;
        RECT  0.740 1.015 0.970 2.900 ;
        RECT  0.275 2.380 0.505 3.430 ;
    END
END AO221D2BWP7T

MACRO AO222D0BWP7T
    CLASS CORE ;
    FOREIGN AO222D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 0.575 6.020 2.805 ;
        RECT  5.695 0.575 5.740 0.915 ;
        RECT  5.695 2.465 5.740 2.805 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.210 4.900 2.150 ;
        RECT  4.500 1.730 4.620 2.150 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 1.210 3.785 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.450 1.155 2.495 1.385 ;
        RECT  0.140 1.155 0.450 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.150 ;
        RECT  2.615 1.805 2.940 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.105 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 1.650 1.030 1.990 ;
        RECT  0.700 1.650 1.010 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.090 -0.235 6.160 0.235 ;
        RECT  4.710 -0.235 5.090 0.820 ;
        RECT  2.215 -0.235 4.710 0.235 ;
        RECT  1.875 -0.235 2.215 0.465 ;
        RECT  0.000 -0.235 1.875 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.420 3.685 6.160 4.155 ;
        RECT  5.080 3.455 5.420 4.155 ;
        RECT  3.960 3.685 5.080 4.155 ;
        RECT  3.620 3.455 3.960 4.155 ;
        RECT  0.000 3.685 3.620 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.140 1.115 5.370 2.610 ;
        RECT  4.245 2.380 5.140 2.610 ;
        RECT  3.090 2.840 4.720 3.070 ;
        RECT  4.015 0.595 4.245 2.610 ;
        RECT  3.410 0.595 4.015 0.825 ;
        RECT  1.805 2.380 4.015 2.610 ;
        RECT  3.175 0.595 3.410 0.925 ;
        RECT  1.120 0.695 3.175 0.925 ;
        RECT  2.860 2.840 3.090 3.445 ;
        RECT  0.520 3.215 2.860 3.445 ;
        RECT  1.575 2.380 1.805 2.970 ;
        RECT  0.890 0.595 1.120 0.925 ;
        RECT  0.610 0.595 0.890 0.825 ;
        RECT  0.180 2.980 0.520 3.445 ;
    END
END AO222D0BWP7T

MACRO AO222D1BWP7T
    CLASS CORE ;
    FOREIGN AO222D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.240 0.495 6.580 3.325 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.670 5.460 2.710 ;
        RECT  4.960 1.670 5.180 2.010 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.730 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.660 2.150 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.755 -0.235 6.720 0.235 ;
        RECT  5.375 -0.235 5.755 0.935 ;
        RECT  3.275 -0.235 5.375 0.235 ;
        RECT  2.895 -0.235 3.275 0.935 ;
        RECT  0.465 -0.235 2.895 0.235 ;
        RECT  0.235 -0.235 0.465 1.245 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 3.685 6.720 4.155 ;
        RECT  5.380 3.025 5.760 4.155 ;
        RECT  4.230 3.685 5.380 4.155 ;
        RECT  3.850 3.085 4.230 4.155 ;
        RECT  0.000 3.685 3.850 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.765 1.190 5.995 2.000 ;
        RECT  4.960 1.190 5.765 1.420 ;
        RECT  4.720 0.685 4.960 1.420 ;
        RECT  4.635 2.490 4.865 3.325 ;
        RECT  3.800 0.685 4.720 0.915 ;
        RECT  2.400 2.490 4.635 2.720 ;
        RECT  3.560 0.685 3.800 1.420 ;
        RECT  2.620 1.190 3.560 1.420 ;
        RECT  0.180 3.085 3.460 3.315 ;
        RECT  2.380 0.695 2.620 1.420 ;
        RECT  0.960 0.695 2.380 0.925 ;
        RECT  0.960 2.565 1.240 2.795 ;
        RECT  0.730 0.695 0.960 2.795 ;
    END
END AO222D1BWP7T

MACRO AO222D2BWP7T
    CLASS CORE ;
    FOREIGN AO222D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.325 0.705 6.580 2.725 ;
        RECT  6.300 0.705 6.325 3.405 ;
        RECT  6.040 0.705 6.300 0.935 ;
        RECT  6.095 2.455 6.300 3.405 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.735 5.460 2.150 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.670 4.370 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.705 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.660 2.150 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 -0.235 7.280 0.235 ;
        RECT  6.815 -0.235 7.045 1.285 ;
        RECT  5.680 -0.235 6.815 0.235 ;
        RECT  5.300 -0.235 5.680 0.935 ;
        RECT  3.280 -0.235 5.300 0.235 ;
        RECT  2.900 -0.235 3.280 0.935 ;
        RECT  0.465 -0.235 2.900 0.235 ;
        RECT  0.235 -0.235 0.465 1.270 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 3.685 7.280 4.155 ;
        RECT  6.815 2.245 7.045 4.155 ;
        RECT  5.680 3.685 6.815 4.155 ;
        RECT  5.300 2.500 5.680 4.155 ;
        RECT  4.230 3.685 5.300 4.155 ;
        RECT  3.850 2.950 4.230 4.155 ;
        RECT  0.000 3.685 3.850 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.815 1.190 6.045 1.985 ;
        RECT  4.155 1.190 5.815 1.420 ;
        RECT  4.635 2.485 4.865 3.295 ;
        RECT  2.400 2.485 4.635 2.715 ;
        RECT  3.905 0.495 4.155 1.420 ;
        RECT  2.620 1.190 3.905 1.420 ;
        RECT  0.160 3.085 3.460 3.315 ;
        RECT  2.380 0.695 2.620 1.420 ;
        RECT  0.960 0.695 2.380 0.925 ;
        RECT  0.960 2.565 1.245 2.795 ;
        RECT  0.730 0.695 0.960 2.795 ;
    END
END AO222D2BWP7T

MACRO AO22D0BWP7T
    CLASS CORE ;
    FOREIGN AO22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5747 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 0.540 4.340 3.300 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.050 1.260 3.280 2.340 ;
        RECT  1.090 1.260 3.050 1.540 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.770 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.385 -0.235 4.480 0.235 ;
        RECT  3.045 -0.235 3.385 0.465 ;
        RECT  0.520 -0.235 3.045 0.235 ;
        RECT  0.180 -0.235 0.520 0.825 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.575 3.685 4.480 4.155 ;
        RECT  3.235 3.030 3.575 4.155 ;
        RECT  0.520 3.685 3.235 4.155 ;
        RECT  0.180 3.030 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.530 0.695 3.760 2.800 ;
        RECT  1.720 0.695 3.530 0.925 ;
        RECT  2.135 2.570 3.530 2.800 ;
        RECT  2.745 3.030 2.855 3.260 ;
        RECT  2.515 3.030 2.745 3.455 ;
        RECT  1.230 3.225 2.515 3.455 ;
        RECT  1.795 2.570 2.135 2.995 ;
        RECT  1.490 0.525 1.720 0.925 ;
        RECT  1.000 2.975 1.230 3.455 ;
    END
END AO22D0BWP7T

MACRO AO22D1BWP7T
    CLASS CORE ;
    FOREIGN AO22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 0.495 4.900 3.370 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.715 1.540 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.730 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 1.655 3.780 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.155 -0.235 5.040 0.235 ;
        RECT  3.780 -0.235 4.155 0.860 ;
        RECT  1.960 -0.235 3.780 0.235 ;
        RECT  1.550 -0.235 1.960 0.885 ;
        RECT  0.000 -0.235 1.550 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.090 3.685 5.040 4.155 ;
        RECT  3.845 3.040 4.090 4.155 ;
        RECT  1.275 3.685 3.845 4.155 ;
        RECT  0.895 2.985 1.275 4.155 ;
        RECT  0.000 3.685 0.895 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.045 1.160 4.275 2.745 ;
        RECT  3.245 1.160 4.045 1.390 ;
        RECT  2.355 2.515 4.045 2.745 ;
        RECT  1.865 2.995 3.415 3.225 ;
        RECT  3.015 0.495 3.245 1.390 ;
        RECT  1.240 1.160 3.015 1.390 ;
        RECT  1.635 2.470 1.865 3.225 ;
        RECT  0.465 2.470 1.635 2.700 ;
        RECT  1.005 0.720 1.240 1.390 ;
        RECT  0.240 0.720 1.005 0.950 ;
        RECT  0.235 2.470 0.465 3.280 ;
    END
END AO22D1BWP7T

MACRO AO22D2BWP7T
    CLASS CORE ;
    FOREIGN AO22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.3154 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.645 0.720 4.900 2.625 ;
        RECT  4.620 0.720 4.645 3.380 ;
        RECT  4.360 0.720 4.620 0.950 ;
        RECT  4.415 2.395 4.620 3.380 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.725 1.540 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.695 3.780 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.365 -0.235 5.600 0.235 ;
        RECT  5.135 -0.235 5.365 1.260 ;
        RECT  3.975 -0.235 5.135 0.235 ;
        RECT  3.605 -0.235 3.975 0.895 ;
        RECT  1.930 -0.235 3.605 0.235 ;
        RECT  1.515 -0.235 1.930 0.465 ;
        RECT  0.000 -0.235 1.515 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.365 3.685 5.600 4.155 ;
        RECT  5.135 2.245 5.365 4.155 ;
        RECT  3.980 3.685 5.135 4.155 ;
        RECT  3.600 3.155 3.980 4.155 ;
        RECT  1.260 3.685 3.600 4.155 ;
        RECT  0.880 2.940 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.160 1.200 4.390 2.000 ;
        RECT  3.285 1.200 4.160 1.430 ;
        RECT  3.115 2.385 3.345 3.340 ;
        RECT  3.030 0.710 3.285 1.430 ;
        RECT  1.905 3.110 3.115 3.340 ;
        RECT  2.625 0.710 3.030 0.940 ;
        RECT  2.395 0.710 2.625 2.690 ;
        RECT  0.180 0.710 2.395 0.940 ;
        RECT  1.675 2.480 1.905 3.340 ;
        RECT  0.465 2.480 1.675 2.710 ;
        RECT  0.235 2.480 0.465 3.320 ;
    END
END AO22D2BWP7T

MACRO AO31D0BWP7T
    CLASS CORE ;
    FOREIGN AO31D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5806 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 0.525 4.340 3.125 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.210 1.540 2.190 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.190 2.105 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.510 -0.235 4.480 0.235 ;
        RECT  3.130 -0.235 3.510 0.785 ;
        RECT  0.580 -0.235 3.130 0.235 ;
        RECT  0.200 -0.235 0.580 0.825 ;
        RECT  0.000 -0.235 0.200 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 3.685 4.480 4.155 ;
        RECT  3.185 2.905 3.565 4.155 ;
        RECT  0.000 3.685 3.185 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.525 1.060 3.755 2.665 ;
        RECT  2.565 1.060 3.525 1.290 ;
        RECT  1.990 2.435 3.525 2.665 ;
        RECT  2.525 2.920 2.755 3.455 ;
        RECT  2.335 0.545 2.565 1.290 ;
        RECT  1.225 3.225 2.525 3.455 ;
        RECT  1.760 2.435 1.990 2.995 ;
        RECT  0.505 2.435 1.760 2.665 ;
        RECT  0.995 2.920 1.225 3.455 ;
        RECT  0.275 2.435 0.505 3.130 ;
    END
END AO31D0BWP7T

MACRO AO31D1BWP7T
    CLASS CORE ;
    FOREIGN AO31D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1444 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 0.495 4.340 3.380 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 1.210 3.220 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.455 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 0.650 1.540 1.855 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.660 2.245 2.150 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 -0.235 4.480 0.235 ;
        RECT  3.135 -0.235 3.495 0.465 ;
        RECT  0.600 -0.235 3.135 0.235 ;
        RECT  0.220 -0.235 0.600 0.970 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.560 3.685 4.480 4.155 ;
        RECT  3.180 3.155 3.560 4.155 ;
        RECT  0.000 3.685 3.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.520 0.695 3.750 2.715 ;
        RECT  2.590 0.695 3.520 0.925 ;
        RECT  0.525 2.485 3.520 2.715 ;
        RECT  0.960 2.990 2.805 3.220 ;
        RECT  2.360 0.495 2.590 1.305 ;
        RECT  0.295 2.485 0.525 3.295 ;
    END
END AO31D1BWP7T

MACRO AO31D2BWP7T
    CLASS CORE ;
    FOREIGN AO31D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.065 0.585 4.340 2.620 ;
        RECT  4.060 0.585 4.065 3.390 ;
        RECT  3.835 0.585 4.060 0.970 ;
        RECT  3.835 2.385 4.060 3.390 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.680 3.220 2.710 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.490 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 0.650 1.540 1.850 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.130 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 -0.235 5.040 0.235 ;
        RECT  4.575 -0.235 4.805 1.260 ;
        RECT  3.425 -0.235 4.575 0.235 ;
        RECT  3.045 -0.235 3.425 0.785 ;
        RECT  0.555 -0.235 3.045 0.235 ;
        RECT  0.175 -0.235 0.555 0.940 ;
        RECT  0.000 -0.235 0.175 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 3.685 5.040 4.155 ;
        RECT  4.575 2.250 4.805 4.155 ;
        RECT  3.420 3.685 4.575 4.155 ;
        RECT  3.040 3.140 3.420 4.155 ;
        RECT  0.000 3.685 3.040 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.600 1.220 3.830 2.020 ;
        RECT  2.590 1.220 3.600 1.450 ;
        RECT  0.900 3.155 2.680 3.385 ;
        RECT  2.360 0.495 2.590 2.815 ;
        RECT  0.465 2.585 2.360 2.815 ;
        RECT  0.235 2.585 0.465 3.395 ;
    END
END AO31D2BWP7T

MACRO AO32D0BWP7T
    CLASS CORE ;
    FOREIGN AO32D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 0.530 5.460 3.280 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.760 4.340 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.765 3.250 2.710 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.570 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.170 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.400 -0.235 5.600 0.235 ;
        RECT  4.020 -0.235 4.400 0.805 ;
        RECT  0.560 -0.235 4.020 0.235 ;
        RECT  0.175 -0.235 0.560 0.815 ;
        RECT  0.000 -0.235 0.175 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.360 3.685 5.600 4.155 ;
        RECT  4.020 3.455 4.360 4.155 ;
        RECT  0.000 3.685 4.020 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.635 1.170 4.865 1.985 ;
        RECT  2.645 1.170 4.635 1.400 ;
        RECT  3.740 2.565 4.145 2.795 ;
        RECT  3.510 2.565 3.740 3.335 ;
        RECT  2.695 3.105 3.510 3.335 ;
        RECT  2.355 2.910 2.695 3.335 ;
        RECT  2.640 1.170 2.645 2.680 ;
        RECT  2.410 0.525 2.640 2.680 ;
        RECT  1.980 2.450 2.410 2.680 ;
        RECT  1.255 3.105 2.355 3.335 ;
        RECT  1.635 2.450 1.980 2.875 ;
        RECT  0.475 2.450 1.635 2.680 ;
        RECT  0.915 2.910 1.255 3.335 ;
        RECT  0.245 2.450 0.475 3.060 ;
    END
END AO32D0BWP7T

MACRO AO32D1BWP7T
    CLASS CORE ;
    FOREIGN AO32D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 0.485 5.460 3.375 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.825 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.210 3.220 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.735 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.650 2.150 1.900 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.405 -0.235 5.600 0.235 ;
        RECT  4.025 -0.235 4.405 0.465 ;
        RECT  0.550 -0.235 4.025 0.235 ;
        RECT  0.170 -0.235 0.550 0.785 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.645 3.685 5.600 4.155 ;
        RECT  4.415 2.335 4.645 4.155 ;
        RECT  3.400 3.685 4.415 4.155 ;
        RECT  3.060 3.250 3.400 4.155 ;
        RECT  0.000 3.685 3.060 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.655 0.695 4.885 2.020 ;
        RECT  2.615 0.695 4.655 0.925 ;
        RECT  3.835 2.790 4.065 3.455 ;
        RECT  2.825 2.790 3.835 3.020 ;
        RECT  2.560 2.790 2.825 3.210 ;
        RECT  2.385 0.465 2.615 2.420 ;
        RECT  0.870 2.980 2.560 3.210 ;
        RECT  2.240 2.190 2.385 2.420 ;
        RECT  2.000 2.190 2.240 2.650 ;
        RECT  0.465 2.420 2.000 2.650 ;
        RECT  0.235 2.420 0.465 3.385 ;
    END
END AO32D1BWP7T

MACRO AO32D2BWP7T
    CLASS CORE ;
    FOREIGN AO32D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.765 1.165 6.020 2.575 ;
        RECT  5.740 0.465 5.765 3.420 ;
        RECT  5.535 0.465 5.740 1.440 ;
        RECT  5.535 2.345 5.740 3.420 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.680 4.340 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.880 1.680 3.245 2.710 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.700 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.210 1.560 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.155 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 -0.235 6.720 0.235 ;
        RECT  6.255 -0.235 6.485 1.270 ;
        RECT  5.120 -0.235 6.255 0.235 ;
        RECT  4.740 -0.235 5.120 0.785 ;
        RECT  4.145 -0.235 4.740 0.235 ;
        RECT  3.765 -0.235 4.145 0.785 ;
        RECT  0.470 -0.235 3.765 0.235 ;
        RECT  0.240 -0.235 0.470 1.305 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 3.685 6.720 4.155 ;
        RECT  6.255 2.250 6.485 4.155 ;
        RECT  5.045 3.685 6.255 4.155 ;
        RECT  4.815 2.250 5.045 4.155 ;
        RECT  3.445 3.685 4.815 4.155 ;
        RECT  3.105 3.455 3.445 4.155 ;
        RECT  0.000 3.685 3.105 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.955 1.020 5.185 2.010 ;
        RECT  2.620 1.020 4.955 1.260 ;
        RECT  3.920 2.380 4.150 3.190 ;
        RECT  0.845 2.960 3.920 3.190 ;
        RECT  2.390 0.465 2.620 2.610 ;
        RECT  0.470 2.380 2.390 2.610 ;
        RECT  0.240 2.380 0.470 3.385 ;
    END
END AO32D2BWP7T

MACRO AO33D0BWP7T
    CLASS CORE ;
    FOREIGN AO33D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 0.585 5.460 2.750 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.040 1.170 4.340 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.160 3.780 2.150 ;
        RECT  3.375 1.725 3.500 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.730 2.865 2.150 ;
        RECT  2.380 1.210 2.660 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.470 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.535 -0.235 5.600 0.235 ;
        RECT  4.195 -0.235 4.535 0.465 ;
        RECT  0.465 -0.235 4.195 0.235 ;
        RECT  0.235 -0.235 0.465 0.920 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.680 3.685 5.600 4.155 ;
        RECT  4.300 3.455 4.680 4.155 ;
        RECT  3.440 3.685 4.300 4.155 ;
        RECT  3.100 3.455 3.440 4.155 ;
        RECT  0.000 3.685 3.100 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.655 0.700 4.885 2.090 ;
        RECT  0.965 0.700 4.655 0.930 ;
        RECT  2.625 2.490 4.020 2.720 ;
        RECT  2.395 2.490 2.625 3.410 ;
        RECT  1.240 3.180 2.395 3.410 ;
        RECT  1.675 2.380 1.905 2.950 ;
        RECT  0.965 2.380 1.675 2.610 ;
        RECT  0.900 2.840 1.240 3.410 ;
        RECT  0.735 0.700 0.965 2.610 ;
        RECT  0.465 2.380 0.735 2.610 ;
        RECT  0.235 2.380 0.465 3.000 ;
    END
END AO33D0BWP7T

MACRO AO33D1BWP7T
    CLASS CORE ;
    FOREIGN AO33D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.695 0.485 6.020 3.405 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.710 4.900 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.825 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.705 3.220 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.470 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 1.210 1.560 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.145 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 -0.235 6.160 0.235 ;
        RECT  4.695 -0.235 5.075 0.785 ;
        RECT  0.465 -0.235 4.695 0.235 ;
        RECT  0.235 -0.235 0.465 0.915 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.980 3.685 6.160 4.155 ;
        RECT  4.750 2.450 4.980 4.155 ;
        RECT  3.345 3.685 4.750 4.155 ;
        RECT  3.115 2.890 3.345 4.155 ;
        RECT  0.000 3.685 3.115 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.215 1.055 5.445 2.010 ;
        RECT  4.375 1.055 5.215 1.285 ;
        RECT  4.145 0.475 4.375 1.285 ;
        RECT  2.605 0.475 4.145 0.705 ;
        RECT  3.855 2.420 4.085 3.415 ;
        RECT  2.625 2.420 3.855 2.650 ;
        RECT  2.395 2.420 2.625 3.310 ;
        RECT  2.375 0.475 2.605 1.285 ;
        RECT  0.895 3.075 2.395 3.310 ;
        RECT  0.930 0.475 2.375 0.705 ;
        RECT  0.930 2.475 1.985 2.705 ;
        RECT  0.700 0.475 0.930 2.705 ;
        RECT  0.465 2.475 0.700 2.705 ;
        RECT  0.235 2.475 0.465 3.385 ;
    END
END AO33D1BWP7T

MACRO AO33D2BWP7T
    CLASS CORE ;
    FOREIGN AO33D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.3035 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.755 1.200 6.020 2.575 ;
        RECT  5.740 0.465 5.755 3.430 ;
        RECT  5.525 0.465 5.740 1.440 ;
        RECT  5.525 2.345 5.740 3.430 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.660 4.550 2.000 ;
        RECT  4.060 1.660 4.340 2.710 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.830 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.150 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 -0.235 6.720 0.235 ;
        RECT  6.255 -0.235 6.485 1.235 ;
        RECT  5.110 -0.235 6.255 0.235 ;
        RECT  4.730 -0.235 5.110 0.870 ;
        RECT  0.470 -0.235 4.730 0.235 ;
        RECT  0.240 -0.235 0.470 0.940 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 3.685 6.720 4.155 ;
        RECT  6.255 2.250 6.485 4.155 ;
        RECT  4.915 3.685 6.255 4.155 ;
        RECT  4.685 2.245 4.915 4.155 ;
        RECT  3.350 3.685 4.685 4.155 ;
        RECT  3.120 2.880 3.350 4.155 ;
        RECT  0.000 3.685 3.120 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.065 1.100 5.295 2.010 ;
        RECT  4.450 1.100 5.065 1.330 ;
        RECT  4.220 0.530 4.450 1.330 ;
        RECT  2.625 0.530 4.220 0.760 ;
        RECT  3.830 2.975 4.160 3.205 ;
        RECT  3.600 2.410 3.830 3.205 ;
        RECT  2.635 2.410 3.600 2.640 ;
        RECT  2.400 2.410 2.635 3.290 ;
        RECT  2.395 0.530 2.625 1.285 ;
        RECT  0.865 3.060 2.400 3.290 ;
        RECT  0.935 0.530 2.395 0.760 ;
        RECT  0.935 2.515 1.975 2.745 ;
        RECT  0.705 0.530 0.935 2.745 ;
        RECT  0.470 2.515 0.705 2.745 ;
        RECT  0.240 2.515 0.470 3.340 ;
    END
END AO33D2BWP7T

MACRO AOI211D0BWP7T
    CLASS CORE ;
    FOREIGN AOI211D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.8874 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 0.690 3.185 0.920 ;
        RECT  2.380 0.690 2.660 3.145 ;
        RECT  1.240 1.185 2.380 1.415 ;
        RECT  2.100 2.915 2.380 3.145 ;
        RECT  0.900 0.670 1.240 1.415 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.540 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.820 2.150 2.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.210 3.220 2.170 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 -0.235 3.360 0.235 ;
        RECT  1.645 -0.235 1.995 0.860 ;
        RECT  0.550 -0.235 1.645 0.235 ;
        RECT  0.170 -0.235 0.550 0.900 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 3.685 3.360 4.155 ;
        RECT  0.160 2.810 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
END AOI211D0BWP7T

MACRO AOI211D1BWP7T
    CLASS CORE ;
    FOREIGN AOI211D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.7598 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 0.495 3.125 1.305 ;
        RECT  2.660 1.075 2.895 1.305 ;
        RECT  2.380 1.075 2.660 2.855 ;
        RECT  0.960 2.625 2.380 2.855 ;
        RECT  0.960 0.690 1.240 0.920 ;
        RECT  0.730 0.690 0.960 2.855 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.465 2.710 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.210 1.540 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.135 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 1.680 3.220 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 -0.235 3.360 0.235 ;
        RECT  1.605 -0.235 1.985 0.865 ;
        RECT  0.465 -0.235 1.605 0.235 ;
        RECT  0.235 -0.235 0.465 1.235 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 3.685 3.360 4.155 ;
        RECT  0.155 3.155 0.535 4.155 ;
        RECT  0.000 3.685 0.155 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.400 3.085 3.180 3.315 ;
    END
END AOI211D1BWP7T

MACRO AOI211D2BWP7T
    CLASS CORE ;
    FOREIGN AOI211D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0996 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 0.700 6.020 2.660 ;
        RECT  2.855 0.700 5.740 0.980 ;
        RECT  3.480 2.380 5.740 2.660 ;
        RECT  2.595 0.700 2.855 1.130 ;
        RECT  0.900 0.900 2.595 1.130 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 1.625 2.100 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 1.480 2.840 2.660 ;
        RECT  0.705 2.380 2.610 2.660 ;
        RECT  0.475 1.615 0.705 2.660 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.265 1.260 5.495 1.980 ;
        RECT  3.575 1.260 5.265 1.540 ;
        RECT  3.345 1.260 3.575 1.995 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 1.780 4.950 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 -0.235 6.160 0.235 ;
        RECT  5.640 -0.235 5.980 0.465 ;
        RECT  3.440 -0.235 5.640 0.235 ;
        RECT  3.100 -0.235 3.440 0.465 ;
        RECT  1.990 -0.235 3.100 0.235 ;
        RECT  1.610 -0.235 1.990 0.670 ;
        RECT  0.550 -0.235 1.610 0.235 ;
        RECT  0.170 -0.235 0.550 0.925 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 3.685 6.160 4.155 ;
        RECT  1.440 3.360 1.780 4.155 ;
        RECT  0.000 3.685 1.440 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.180 2.890 5.980 3.120 ;
    END
END AOI211D2BWP7T

MACRO AOI211XD0BWP7T
    CLASS CORE ;
    FOREIGN AOI211XD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2635 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 0.815 3.180 1.045 ;
        RECT  2.380 0.675 2.660 2.995 ;
        RECT  1.200 0.675 2.380 0.905 ;
        RECT  2.110 2.765 2.380 2.995 ;
        RECT  0.940 0.675 1.200 1.125 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.620 0.465 2.710 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 1.625 1.540 2.710 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.105 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.625 3.220 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 -0.235 3.360 0.235 ;
        RECT  0.160 -0.235 0.540 1.045 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 3.685 3.360 4.155 ;
        RECT  0.160 3.045 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.385 3.225 3.180 3.455 ;
    END
END AOI211XD0BWP7T

MACRO AOI211XD1BWP7T
    CLASS CORE ;
    FOREIGN AOI211XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 0.700 6.580 2.660 ;
        RECT  2.065 0.700 6.300 0.980 ;
        RECT  3.860 2.380 6.300 2.660 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 1.770 2.235 2.100 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 1.260 3.185 1.960 ;
        RECT  0.705 1.260 2.955 1.540 ;
        RECT  0.475 1.260 0.705 2.025 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.260 5.970 1.965 ;
        RECT  3.905 1.260 5.740 1.540 ;
        RECT  3.675 1.260 3.905 1.960 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.570 1.770 5.510 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.620 -0.235 6.720 0.235 ;
        RECT  3.280 -0.235 3.620 0.465 ;
        RECT  1.605 -0.235 3.280 0.235 ;
        RECT  1.225 -0.235 1.605 0.950 ;
        RECT  0.000 -0.235 1.225 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 3.685 6.720 4.155 ;
        RECT  1.660 3.450 2.000 4.155 ;
        RECT  0.000 3.685 1.660 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.425 2.990 6.540 3.220 ;
        RECT  3.195 2.390 3.425 3.220 ;
        RECT  0.180 2.990 3.195 3.220 ;
        RECT  0.900 2.490 2.760 2.720 ;
    END
END AOI211XD1BWP7T

MACRO AOI211XD2BWP7T
    CLASS CORE ;
    FOREIGN AOI211XD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.1978 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.380 2.535 11.930 2.765 ;
        RECT  10.080 0.990 10.420 1.385 ;
        RECT  9.380 1.155 10.080 1.385 ;
        RECT  9.100 1.155 9.380 2.765 ;
        RECT  6.645 1.155 9.100 1.385 ;
        RECT  7.000 2.535 9.100 2.765 ;
        RECT  6.415 0.700 6.645 1.385 ;
        RECT  1.000 0.700 6.415 0.980 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.715 3.810 2.150 ;
        RECT  1.590 1.715 2.940 1.945 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.800 1.675 5.860 2.100 ;
        RECT  4.570 1.255 4.800 2.100 ;
        RECT  0.805 1.255 4.570 1.485 ;
        RECT  0.565 1.255 0.805 1.990 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.190 1.695 8.620 1.925 ;
        RECT  6.250 1.695 7.190 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.290 1.695 12.230 2.100 ;
        RECT  9.810 1.695 11.290 1.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.905 -0.235 12.880 0.235 ;
        RECT  8.515 -0.235 8.905 0.465 ;
        RECT  5.240 -0.235 8.515 0.235 ;
        RECT  4.865 -0.235 5.240 0.465 ;
        RECT  3.625 -0.235 4.865 0.235 ;
        RECT  3.275 -0.235 3.625 0.470 ;
        RECT  0.640 -0.235 3.275 0.235 ;
        RECT  0.260 -0.235 0.640 0.930 ;
        RECT  0.000 -0.235 0.260 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.630 3.685 12.880 4.155 ;
        RECT  3.270 3.455 3.630 4.155 ;
        RECT  2.130 3.685 3.270 4.155 ;
        RECT  1.750 3.455 2.130 4.155 ;
        RECT  0.000 3.685 1.750 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.565 2.995 12.625 3.225 ;
        RECT  10.800 0.495 11.140 1.200 ;
        RECT  9.620 0.495 10.800 0.725 ;
        RECT  9.355 0.495 9.620 0.925 ;
        RECT  7.780 0.695 9.355 0.925 ;
        RECT  1.000 2.515 5.820 2.745 ;
        RECT  0.335 2.380 0.565 3.225 ;
    END
END AOI211XD2BWP7T

MACRO AOI21D0BWP7T
    CLASS CORE ;
    FOREIGN AOI21D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6458 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 0.595 1.875 0.825 ;
        RECT  0.980 2.505 1.250 2.735 ;
        RECT  0.700 0.595 0.980 2.735 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.655 2.660 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.575 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.540 -0.235 2.800 0.235 ;
        RECT  2.310 -0.235 2.540 0.850 ;
        RECT  0.470 -0.235 2.310 0.235 ;
        RECT  0.240 -0.235 0.470 0.850 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.640 3.685 2.800 4.155 ;
        RECT  2.270 3.455 2.640 4.155 ;
        RECT  0.000 3.685 2.270 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.690 2.450 1.920 3.210 ;
        RECT  0.470 2.980 1.690 3.210 ;
        RECT  0.240 2.460 0.470 3.210 ;
    END
END AOI21D0BWP7T

MACRO AOI21D1BWP7T
    CLASS CORE ;
    FOREIGN AOI21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.6998 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.535 0.495 2.765 1.345 ;
        RECT  0.980 1.115 2.535 1.345 ;
        RECT  1.095 2.150 1.325 2.895 ;
        RECT  0.980 2.150 1.095 2.380 ;
        RECT  0.700 0.615 0.980 2.380 ;
        RECT  0.320 0.615 0.700 0.845 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.665 3.220 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.645 2.120 2.710 ;
        RECT  1.570 1.645 1.820 1.875 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 -0.235 3.360 0.235 ;
        RECT  1.745 -0.235 2.125 0.825 ;
        RECT  0.000 -0.235 1.745 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 3.685 3.360 4.155 ;
        RECT  2.525 2.455 2.770 4.155 ;
        RECT  0.000 3.685 2.525 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.605 3.225 2.100 3.455 ;
        RECT  0.375 2.595 0.605 3.455 ;
    END
END AOI21D1BWP7T

MACRO AOI21D2BWP7T
    CLASS CORE ;
    FOREIGN AOI21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 2.380 4.150 2.660 ;
        RECT  1.995 0.700 3.420 0.980 ;
        RECT  2.265 2.330 2.550 2.660 ;
        RECT  1.995 2.330 2.265 2.560 ;
        RECT  1.765 0.700 1.995 2.560 ;
        RECT  0.905 0.700 1.765 0.980 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.740 1.305 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.370 1.260 4.600 1.990 ;
        RECT  2.455 1.260 4.370 1.540 ;
        RECT  2.225 1.260 2.455 1.980 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 1.770 3.830 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 -0.235 5.040 0.235 ;
        RECT  4.500 -0.235 4.880 0.960 ;
        RECT  2.005 -0.235 4.500 0.235 ;
        RECT  1.665 -0.235 2.005 0.465 ;
        RECT  0.550 -0.235 1.665 0.235 ;
        RECT  0.170 -0.235 0.550 1.205 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 3.685 5.040 4.155 ;
        RECT  0.885 3.250 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.575 2.350 4.805 3.175 ;
        RECT  1.900 2.945 4.575 3.175 ;
        RECT  1.615 2.790 1.900 3.175 ;
        RECT  0.185 2.790 1.615 3.020 ;
    END
END AOI21D2BWP7T

MACRO AOI221D0BWP7T
    CLASS CORE ;
    FOREIGN AOI221D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.0889 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.670 0.565 3.900 0.980 ;
        RECT  1.590 0.700 3.670 0.980 ;
        RECT  2.480 2.380 2.710 2.920 ;
        RECT  1.590 2.380 2.480 2.660 ;
        RECT  1.560 0.700 1.590 2.660 ;
        RECT  1.360 0.625 1.560 2.660 ;
        RECT  0.945 0.625 1.360 0.855 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.795 1.250 4.025 2.195 ;
        RECT  1.865 1.250 3.795 1.540 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.780 1.120 2.150 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.770 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 3.300 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 -0.235 4.480 0.235 ;
        RECT  2.145 -0.235 2.485 0.465 ;
        RECT  0.560 -0.235 2.145 0.235 ;
        RECT  0.180 -0.235 0.560 0.855 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.560 3.685 4.480 4.155 ;
        RECT  0.180 3.040 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.015 2.570 4.245 3.380 ;
        RECT  1.205 3.150 4.015 3.380 ;
        RECT  0.975 2.965 1.205 3.380 ;
    END
END AOI221D0BWP7T

MACRO AOI221D1BWP7T
    CLASS CORE ;
    FOREIGN AOI221D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.7598 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 0.495 4.900 2.905 ;
        RECT  3.830 0.745 4.575 0.975 ;
        RECT  3.800 2.675 4.575 2.905 ;
        RECT  3.600 0.745 3.830 1.305 ;
        RECT  1.190 1.075 3.600 1.305 ;
        RECT  0.960 0.495 1.190 1.305 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.455 2.150 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.730 2.660 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 1.540 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.735 3.780 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.345 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.370 -0.235 5.040 0.235 ;
        RECT  3.130 -0.235 3.370 0.835 ;
        RECT  2.685 -0.235 3.130 0.235 ;
        RECT  2.340 -0.235 2.685 0.835 ;
        RECT  0.550 -0.235 2.340 0.235 ;
        RECT  0.170 -0.235 0.550 0.880 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 3.685 5.040 4.155 ;
        RECT  0.240 2.470 0.470 4.155 ;
        RECT  0.000 3.685 0.240 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.365 3.155 4.860 3.385 ;
        RECT  3.135 2.675 3.365 3.385 ;
        RECT  1.625 2.675 3.135 2.905 ;
        RECT  1.195 3.155 2.685 3.385 ;
        RECT  0.955 2.490 1.195 3.385 ;
    END
END AOI221D1BWP7T

MACRO AOI221D2BWP7T
    CLASS CORE ;
    FOREIGN AOI221D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 4.9390 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.495 2.350 8.725 3.415 ;
        RECT  8.265 0.495 8.495 1.305 ;
        RECT  5.460 2.675 8.495 2.905 ;
        RECT  5.460 0.695 8.265 0.925 ;
        RECT  5.180 0.695 5.460 2.905 ;
        RECT  4.825 0.695 5.180 0.925 ;
        RECT  4.595 0.495 4.825 1.305 ;
        RECT  1.985 0.695 4.595 0.925 ;
        RECT  1.755 0.495 1.985 1.320 ;
        RECT  0.465 1.090 1.755 1.320 ;
        RECT  0.235 0.495 0.465 1.320 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.600 0.980 2.710 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.780 1.795 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.355 1.635 4.585 2.410 ;
        RECT  2.225 2.180 4.355 2.410 ;
        RECT  1.995 1.680 2.225 2.410 ;
        RECT  1.260 1.680 1.995 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.420 1.210 7.700 1.590 ;
        RECT  6.610 1.210 7.420 1.885 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.650 8.265 2.420 ;
        RECT  6.020 2.180 7.980 2.420 ;
        RECT  5.740 1.590 6.020 2.420 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.210 -0.235 8.960 0.235 ;
        RECT  6.800 -0.235 7.210 0.465 ;
        RECT  3.530 -0.235 6.800 0.235 ;
        RECT  3.160 -0.235 3.530 0.465 ;
        RECT  1.310 -0.235 3.160 0.235 ;
        RECT  0.925 -0.235 1.310 0.790 ;
        RECT  0.000 -0.235 0.925 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 3.685 8.960 4.155 ;
        RECT  0.925 3.430 1.280 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.420 3.155 7.900 3.385 ;
        RECT  2.040 2.675 4.920 2.905 ;
        RECT  1.800 2.675 2.040 3.170 ;
        RECT  0.465 2.940 1.800 3.170 ;
        RECT  0.235 2.440 0.465 3.415 ;
    END
END AOI221D2BWP7T

MACRO AOI222D0BWP7T
    CLASS CORE ;
    FOREIGN AOI222D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.8849 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.020 0.625 4.360 0.860 ;
        RECT  3.835 0.625 4.020 0.950 ;
        RECT  2.030 0.720 3.835 0.950 ;
        RECT  0.980 2.465 3.480 2.695 ;
        RECT  1.840 0.630 2.030 0.950 ;
        RECT  0.980 0.630 1.840 0.860 ;
        RECT  0.700 0.630 0.980 2.695 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.210 1.540 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 1.180 4.900 2.175 ;
        RECT  2.480 1.180 4.575 1.410 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.810 1.210 2.145 2.160 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.225 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.640 4.340 2.710 ;
        RECT  3.620 1.640 4.060 1.870 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.100 -0.235 5.040 0.235 ;
        RECT  2.750 -0.235 3.100 0.465 ;
        RECT  0.470 -0.235 2.750 0.235 ;
        RECT  0.240 -0.235 0.470 0.860 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.170 3.685 5.040 4.155 ;
        RECT  0.830 3.415 1.170 4.155 ;
        RECT  0.000 3.685 0.830 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.575 2.495 4.805 3.170 ;
        RECT  0.465 2.940 4.575 3.170 ;
        RECT  0.235 2.490 0.465 3.170 ;
    END
END AOI222D0BWP7T

MACRO AOI222D1BWP7T
    CLASS CORE ;
    FOREIGN AOI222D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8498 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 0.465 5.365 1.280 ;
        RECT  4.900 1.030 5.135 1.280 ;
        RECT  4.620 1.030 4.900 2.820 ;
        RECT  3.140 1.030 4.620 1.260 ;
        RECT  4.415 2.480 4.620 2.820 ;
        RECT  2.910 0.685 3.140 1.260 ;
        RECT  1.600 0.685 2.910 0.915 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.455 2.150 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.705 1.430 2.150 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.735 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.120 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.735 4.340 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.680 5.460 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.815 -0.235 5.600 0.235 ;
        RECT  3.435 -0.235 3.815 0.785 ;
        RECT  0.545 -0.235 3.435 0.235 ;
        RECT  0.160 -0.235 0.545 0.910 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.240 3.685 5.600 4.155 ;
        RECT  0.900 2.925 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.350 3.170 5.420 3.400 ;
        RECT  1.915 2.410 3.410 2.640 ;
        RECT  1.685 2.410 1.915 3.350 ;
        RECT  0.465 2.410 1.685 2.640 ;
        RECT  0.235 2.410 0.465 3.350 ;
    END
END AOI222D1BWP7T

MACRO AOI222D2BWP7T
    CLASS CORE ;
    FOREIGN AOI222D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.6955 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.830 1.140 9.940 2.905 ;
        RECT  9.660 1.140 9.830 3.430 ;
        RECT  9.305 1.140 9.660 1.370 ;
        RECT  9.600 2.675 9.660 3.430 ;
        RECT  6.665 2.675 9.600 2.905 ;
        RECT  9.065 0.560 9.305 1.370 ;
        RECT  7.575 0.560 9.065 0.790 ;
        RECT  7.345 0.560 7.575 1.290 ;
        RECT  5.555 1.060 7.345 1.290 ;
        RECT  5.325 0.570 5.555 1.290 ;
        RECT  3.815 0.570 5.325 0.800 ;
        RECT  3.575 0.570 3.815 1.290 ;
        RECT  2.625 1.060 3.575 1.290 ;
        RECT  2.395 0.570 2.625 1.290 ;
        RECT  1.645 0.570 2.395 0.800 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.535 2.910 2.410 ;
        RECT  0.470 2.180 2.680 2.410 ;
        RECT  0.140 1.210 0.470 2.410 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 2.165 1.930 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.640 1.615 6.020 2.420 ;
        RECT  3.790 2.180 5.640 2.420 ;
        RECT  3.500 1.565 3.790 2.420 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 5.095 1.855 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.635 9.390 2.410 ;
        RECT  7.140 2.180 9.100 2.410 ;
        RECT  6.860 1.525 7.140 2.410 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.870 1.210 8.820 1.875 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.790 -0.235 10.080 0.235 ;
        RECT  9.560 -0.235 9.790 0.840 ;
        RECT  7.035 -0.235 9.560 0.235 ;
        RECT  6.655 -0.235 7.035 0.785 ;
        RECT  6.190 -0.235 6.655 0.235 ;
        RECT  5.850 -0.235 6.190 0.785 ;
        RECT  3.295 -0.235 5.850 0.235 ;
        RECT  2.915 -0.235 3.295 0.695 ;
        RECT  0.565 -0.235 2.915 0.235 ;
        RECT  0.185 -0.235 0.565 0.910 ;
        RECT  0.000 -0.235 0.185 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.725 3.685 10.080 4.155 ;
        RECT  2.345 3.155 2.725 4.155 ;
        RECT  1.280 3.685 2.345 4.155 ;
        RECT  0.900 3.155 1.280 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.805 3.155 9.165 3.385 ;
        RECT  3.370 2.675 6.305 2.905 ;
        RECT  3.140 2.675 3.370 3.430 ;
        RECT  1.930 2.675 3.140 2.905 ;
        RECT  1.700 2.675 1.930 3.430 ;
        RECT  0.550 2.675 1.700 2.905 ;
        RECT  0.205 2.675 0.550 3.430 ;
    END
END AOI222D2BWP7T

MACRO AOI22D0BWP7T
    CLASS CORE ;
    FOREIGN AOI22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6674 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.930 0.465 1.855 0.695 ;
        RECT  0.980 2.880 1.845 3.110 ;
        RECT  0.930 1.535 0.980 3.110 ;
        RECT  0.700 0.465 0.930 3.110 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.455 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 2.465 3.195 2.695 ;
        RECT  2.380 1.040 2.660 2.695 ;
        RECT  1.160 1.040 2.380 1.270 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.210 3.220 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.205 -0.235 3.360 0.235 ;
        RECT  2.825 -0.235 3.205 0.710 ;
        RECT  0.465 -0.235 2.825 0.235 ;
        RECT  0.235 -0.235 0.465 0.765 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 3.685 3.360 4.155 ;
        RECT  2.895 3.055 3.125 4.155 ;
        RECT  0.465 3.685 2.895 4.155 ;
        RECT  0.235 2.975 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
END AOI22D0BWP7T

MACRO AOI22D1BWP7T
    CLASS CORE ;
    FOREIGN AOI22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.0212 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 0.490 3.780 2.790 ;
        RECT  0.200 0.700 3.455 0.980 ;
        RECT  2.590 2.560 3.455 2.790 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.705 1.540 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.745 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.185 -0.235 3.920 0.235 ;
        RECT  1.845 -0.235 2.185 0.465 ;
        RECT  0.000 -0.235 1.845 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 3.685 3.920 4.155 ;
        RECT  0.960 2.930 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.005 3.115 3.740 3.345 ;
        RECT  1.775 2.380 2.005 3.345 ;
        RECT  0.485 2.380 1.775 2.610 ;
        RECT  0.255 2.380 0.485 3.380 ;
    END
END AOI22D1BWP7T

MACRO AOI22D2BWP7T
    CLASS CORE ;
    FOREIGN AOI22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.6270 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 0.715 6.580 2.810 ;
        RECT  1.680 0.715 6.300 0.945 ;
        RECT  3.940 2.580 6.300 2.810 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.210 3.220 2.150 ;
        RECT  0.980 1.210 2.855 1.440 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.745 2.250 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.190 6.020 2.150 ;
        RECT  3.780 1.190 5.740 1.420 ;
        RECT  3.500 1.190 3.780 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.415 1.735 5.460 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.445 -0.235 6.720 0.235 ;
        RECT  6.040 -0.235 6.445 0.465 ;
        RECT  3.540 -0.235 6.040 0.235 ;
        RECT  3.110 -0.235 3.540 0.465 ;
        RECT  0.470 -0.235 3.110 0.235 ;
        RECT  0.240 -0.235 0.470 1.250 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.775 3.685 6.720 4.155 ;
        RECT  2.395 2.930 2.775 4.155 ;
        RECT  1.295 3.685 2.395 4.155 ;
        RECT  0.915 2.930 1.295 4.155 ;
        RECT  0.000 3.685 0.915 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.465 3.155 6.480 3.385 ;
        RECT  3.235 2.470 3.465 3.385 ;
        RECT  1.965 2.470 3.235 2.700 ;
        RECT  1.735 2.470 1.965 3.280 ;
        RECT  0.470 2.470 1.735 2.700 ;
        RECT  0.240 2.470 0.470 3.365 ;
    END
END AOI22D2BWP7T

MACRO AOI31D0BWP7T
    CLASS CORE ;
    FOREIGN AOI31D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9921 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.630 2.660 2.705 ;
        RECT  2.085 0.630 2.380 0.860 ;
        RECT  0.180 2.475 2.380 2.705 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.900 1.210 3.220 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.165 0.650 1.540 1.605 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.105 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.235 3.360 0.235 ;
        RECT  2.895 -0.235 3.125 0.885 ;
        RECT  0.465 -0.235 2.895 0.235 ;
        RECT  0.235 -0.235 0.465 0.895 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 3.685 3.360 4.155 ;
        RECT  2.895 2.440 3.125 4.155 ;
        RECT  0.000 3.685 2.895 4.155 ;
        END
    END VDD
END AOI31D0BWP7T

MACRO AOI31D1BWP7T
    CLASS CORE ;
    FOREIGN AOI31D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.1944 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 0.650 2.740 0.880 ;
        RECT  1.820 0.650 2.100 2.660 ;
        RECT  0.525 2.380 1.820 2.660 ;
        RECT  0.295 2.380 0.525 3.350 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.255 1.210 3.780 1.590 ;
        RECT  2.940 1.210 3.255 1.915 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 0.640 1.540 1.855 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 1.200 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.570 -0.235 3.920 0.235 ;
        RECT  3.190 -0.235 3.570 0.895 ;
        RECT  0.600 -0.235 3.190 0.235 ;
        RECT  0.220 -0.235 0.600 0.900 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 3.685 3.920 4.155 ;
        RECT  3.260 2.250 3.495 4.155 ;
        RECT  0.000 3.685 3.260 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.515 2.410 2.745 3.405 ;
        RECT  0.960 2.890 2.515 3.120 ;
    END
END AOI31D1BWP7T

MACRO AOI31D2BWP7T
    CLASS CORE ;
    FOREIGN AOI31D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.1906 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 0.700 6.580 2.995 ;
        RECT  0.930 0.700 6.300 0.980 ;
        RECT  2.370 2.765 6.300 2.995 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8280 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.705 1.540 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.8064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.365 6.060 2.535 ;
        RECT  2.435 2.305 5.740 2.535 ;
        RECT  2.195 1.770 2.435 2.535 ;
        RECT  1.820 1.770 2.195 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.7785 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 1.260 5.440 1.685 ;
        RECT  3.540 1.260 5.100 1.540 ;
        RECT  3.200 1.260 3.540 1.615 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.7785 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.845 4.280 2.075 ;
        RECT  2.700 1.260 2.930 2.075 ;
        RECT  1.770 1.260 2.700 1.540 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.540 -0.235 6.720 0.235 ;
        RECT  6.200 -0.235 6.540 0.465 ;
        RECT  2.120 -0.235 6.200 0.235 ;
        RECT  1.775 -0.235 2.120 0.470 ;
        RECT  0.560 -0.235 1.775 0.235 ;
        RECT  0.180 -0.235 0.560 0.915 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.295 3.685 6.720 4.155 ;
        RECT  0.915 3.035 1.295 4.155 ;
        RECT  0.000 3.685 0.915 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.935 3.225 6.540 3.455 ;
        RECT  1.705 2.495 1.935 3.455 ;
        RECT  0.490 2.495 1.705 2.725 ;
        RECT  0.260 2.495 0.490 3.415 ;
    END
END AOI31D2BWP7T

MACRO AOI32D0BWP7T
    CLASS CORE ;
    FOREIGN AOI32D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.705 2.660 2.610 ;
        RECT  2.010 2.380 2.380 2.610 ;
        RECT  1.670 2.380 2.010 2.805 ;
        RECT  0.510 2.380 1.670 2.610 ;
        RECT  0.280 2.380 0.510 2.990 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 4.340 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.700 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.145 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.130 -0.235 4.480 0.235 ;
        RECT  3.900 -0.235 4.130 1.060 ;
        RECT  0.515 -0.235 3.900 0.235 ;
        RECT  0.275 -0.235 0.515 1.070 ;
        RECT  0.000 -0.235 0.275 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 3.685 4.480 4.155 ;
        RECT  3.185 3.300 3.525 4.155 ;
        RECT  0.000 3.685 3.185 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.745 2.840 4.300 3.070 ;
        RECT  2.405 2.840 2.745 3.265 ;
        RECT  1.290 3.035 2.405 3.265 ;
        RECT  0.950 2.840 1.290 3.265 ;
    END
END AOI32D0BWP7T

MACRO AOI32D1BWP7T
    CLASS CORE ;
    FOREIGN AOI32D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.4051 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 0.465 2.705 1.290 ;
        RECT  0.980 0.700 2.475 0.980 ;
        RECT  0.980 2.550 2.020 2.790 ;
        RECT  0.700 0.700 0.980 2.790 ;
        RECT  0.525 2.500 0.700 2.790 ;
        RECT  0.295 2.500 0.525 3.310 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.730 4.340 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.715 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 -0.235 4.480 0.235 ;
        RECT  3.910 -0.235 4.140 1.280 ;
        RECT  0.470 -0.235 3.910 0.235 ;
        RECT  0.240 -0.235 0.470 0.925 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 3.685 4.480 4.155 ;
        RECT  3.120 3.065 3.500 4.155 ;
        RECT  0.000 3.685 3.120 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.910 2.520 4.140 3.400 ;
        RECT  2.700 2.520 3.910 2.750 ;
        RECT  2.470 2.520 2.700 3.385 ;
        RECT  0.960 3.155 2.470 3.385 ;
    END
END AOI32D1BWP7T

MACRO AOI32D2BWP7T
    CLASS CORE ;
    FOREIGN AOI32D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.5015 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 0.660 8.260 2.940 ;
        RECT  7.760 0.660 8.030 0.900 ;
        RECT  3.825 2.710 8.030 2.940 ;
        RECT  3.780 0.700 4.075 0.930 ;
        RECT  3.780 1.890 3.825 2.940 ;
        RECT  3.585 0.700 3.780 2.940 ;
        RECT  3.500 0.700 3.585 2.150 ;
        RECT  1.510 0.700 3.500 0.930 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.645 1.210 2.875 1.980 ;
        RECT  0.455 1.210 2.645 1.470 ;
        RECT  0.140 1.210 0.455 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 1.700 2.110 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.610 1.210 6.580 1.840 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.835 0.700 7.065 1.885 ;
        RECT  4.955 0.700 6.835 0.980 ;
        RECT  4.725 0.700 4.955 1.750 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.420 1.390 7.735 2.355 ;
        RECT  4.340 2.125 7.420 2.355 ;
        RECT  4.055 1.770 4.340 2.355 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.115 -0.235 8.400 0.235 ;
        RECT  5.775 -0.235 6.115 0.465 ;
        RECT  3.260 -0.235 5.775 0.235 ;
        RECT  2.910 -0.235 3.260 0.465 ;
        RECT  0.550 -0.235 2.910 0.235 ;
        RECT  0.170 -0.235 0.550 0.910 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.705 3.685 8.400 4.155 ;
        RECT  2.325 3.035 2.705 4.155 ;
        RECT  1.265 3.685 2.325 4.155 ;
        RECT  0.885 3.040 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.355 3.225 8.165 3.455 ;
        RECT  3.125 2.510 3.355 3.455 ;
        RECT  1.915 2.510 3.125 2.740 ;
        RECT  1.685 2.510 1.915 3.320 ;
        RECT  0.470 2.510 1.685 2.740 ;
        RECT  0.240 2.510 0.470 3.320 ;
    END
END AOI32D2BWP7T

MACRO AOI33D0BWP7T
    CLASS CORE ;
    FOREIGN AOI33D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1590 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 0.585 2.655 0.815 ;
        RECT  1.625 2.400 1.965 2.995 ;
        RECT  0.980 2.400 1.625 2.630 ;
        RECT  0.700 0.585 0.980 2.630 ;
        RECT  0.465 2.400 0.700 2.630 ;
        RECT  0.235 2.400 0.465 3.185 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.720 4.920 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.180 3.780 2.190 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 1.210 3.220 2.190 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.710 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.765 -0.235 5.040 0.235 ;
        RECT  4.385 -0.235 4.765 0.805 ;
        RECT  0.465 -0.235 4.385 0.235 ;
        RECT  0.235 -0.235 0.465 0.855 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 3.685 5.040 4.155 ;
        RECT  4.575 2.835 4.805 4.155 ;
        RECT  3.365 3.685 4.575 4.155 ;
        RECT  3.135 2.905 3.365 4.155 ;
        RECT  0.000 3.685 3.135 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.855 2.435 4.085 3.185 ;
        RECT  2.645 2.435 3.855 2.665 ;
        RECT  2.415 2.435 2.645 3.455 ;
        RECT  1.190 3.225 2.415 3.455 ;
        RECT  0.960 2.865 1.190 3.455 ;
    END
END AOI33D0BWP7T

MACRO AOI33D1BWP7T
    CLASS CORE ;
    FOREIGN AOI33D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.1780 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 0.670 2.570 0.900 ;
        RECT  0.980 2.530 1.970 2.760 ;
        RECT  0.700 0.670 0.980 2.760 ;
        RECT  0.465 2.530 0.700 2.760 ;
        RECT  0.235 2.530 0.465 3.340 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.705 4.900 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.210 3.220 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.165 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.685 -0.235 5.040 0.235 ;
        RECT  4.455 -0.235 4.685 1.310 ;
        RECT  0.465 -0.235 4.455 0.235 ;
        RECT  0.235 -0.235 0.465 0.980 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 3.685 5.040 4.155 ;
        RECT  4.575 2.455 4.805 4.155 ;
        RECT  3.365 3.685 4.575 4.155 ;
        RECT  3.135 2.950 3.365 4.155 ;
        RECT  0.000 3.685 3.135 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.855 2.455 4.085 3.450 ;
        RECT  2.645 2.455 3.855 2.685 ;
        RECT  2.415 2.455 2.645 3.325 ;
        RECT  0.900 3.095 2.415 3.325 ;
    END
END AOI33D1BWP7T

MACRO AOI33D2BWP7T
    CLASS CORE ;
    FOREIGN AOI33D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.4318 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.175 0.625 9.405 2.995 ;
        RECT  8.975 0.625 9.175 0.905 ;
        RECT  5.280 2.765 9.175 2.995 ;
        RECT  5.200 0.665 5.430 1.185 ;
        RECT  5.050 2.330 5.280 2.995 ;
        RECT  4.900 0.955 5.200 1.185 ;
        RECT  4.900 2.330 5.050 2.560 ;
        RECT  4.620 0.955 4.900 2.560 ;
        RECT  4.270 0.955 4.620 1.185 ;
        RECT  4.040 0.465 4.270 1.185 ;
        RECT  2.075 0.465 4.040 0.695 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.810 1.770 4.340 2.150 ;
        RECT  3.580 0.925 3.810 2.150 ;
        RECT  0.980 0.925 3.580 1.155 ;
        RECT  0.700 0.925 0.980 1.720 ;
        RECT  0.415 1.490 0.700 1.720 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.490 3.350 1.730 ;
        RECT  2.940 1.490 3.220 2.560 ;
        RECT  1.540 2.330 2.940 2.560 ;
        RECT  1.245 1.620 1.540 2.560 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.820 2.710 2.100 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.305 1.260 7.750 1.540 ;
        RECT  7.075 1.260 7.305 1.965 ;
        RECT  6.810 1.260 7.075 1.540 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.045 0.700 8.275 1.955 ;
        RECT  6.340 0.700 8.045 0.980 ;
        RECT  6.110 0.700 6.340 1.775 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 1.435 8.945 1.775 ;
        RECT  8.540 1.210 8.820 2.535 ;
        RECT  5.770 2.305 8.540 2.535 ;
        RECT  5.540 1.680 5.770 2.535 ;
        RECT  5.225 1.680 5.540 1.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.350 -0.235 9.520 0.235 ;
        RECT  6.990 -0.235 7.350 0.465 ;
        RECT  4.730 -0.235 6.990 0.235 ;
        RECT  4.500 -0.235 4.730 0.725 ;
        RECT  0.465 -0.235 4.500 0.235 ;
        RECT  0.235 -0.235 0.465 0.905 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.120 3.685 9.520 4.155 ;
        RECT  3.780 3.250 4.120 4.155 ;
        RECT  2.680 3.685 3.780 4.155 ;
        RECT  2.340 3.250 2.680 4.155 ;
        RECT  1.240 3.685 2.340 4.155 ;
        RECT  0.895 3.250 1.240 4.155 ;
        RECT  0.000 3.685 0.895 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.785 3.225 9.330 3.455 ;
        RECT  4.555 2.790 4.785 3.455 ;
        RECT  0.465 2.790 4.555 3.020 ;
        RECT  0.235 2.450 0.465 3.435 ;
    END
END AOI33D2BWP7T

MACRO BHDBWP7T
    CLASS CORE ;
    FOREIGN BHDBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNAGATEAREA 0.2133 ;
        ANTENNADIFFAREA 0.4242 ;
        DIRECTION INOUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.730 2.660 3.275 ;
        RECT  2.245 0.730 2.380 0.970 ;
        RECT  0.740 2.150 2.380 2.390 ;
        RECT  2.245 3.035 2.380 3.275 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.340 -0.235 2.800 0.235 ;
        RECT  0.960 -0.235 1.340 0.970 ;
        RECT  0.000 -0.235 0.960 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.340 3.685 2.800 4.155 ;
        RECT  0.960 3.025 1.340 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.470 1.450 1.960 1.690 ;
        RECT  0.230 0.680 0.470 3.190 ;
    END
END BHDBWP7T

MACRO BUFFD0BWP7T
    CLASS CORE ;
    FOREIGN BUFFD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5925 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.685 2.100 3.315 ;
        RECT  1.720 0.685 1.820 0.930 ;
        RECT  1.700 3.075 1.820 3.315 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.235 2.240 0.235 ;
        RECT  0.930 -0.235 1.310 0.910 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 3.685 2.240 4.155 ;
        RECT  0.930 3.065 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.470 2.380 1.560 2.620 ;
        RECT  0.230 0.635 0.470 3.365 ;
    END
END BUFFD0BWP7T

MACRO BUFFD10BWP7T
    CLASS CORE ;
    FOREIGN BUFFD10BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 6.3990 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.450 0.495 9.690 1.390 ;
        RECT  9.450 2.150 9.690 3.365 ;
        RECT  8.230 0.990 9.450 1.390 ;
        RECT  8.230 2.150 9.450 2.550 ;
        RECT  7.990 0.495 8.230 1.390 ;
        RECT  7.990 2.150 8.230 3.365 ;
        RECT  7.450 0.990 7.990 1.390 ;
        RECT  7.450 2.150 7.990 2.550 ;
        RECT  6.790 0.990 7.450 2.550 ;
        RECT  6.550 0.495 6.790 3.365 ;
        RECT  5.990 0.990 6.550 2.550 ;
        RECT  5.350 0.990 5.990 1.390 ;
        RECT  5.350 2.150 5.990 2.550 ;
        RECT  5.110 0.495 5.350 1.390 ;
        RECT  5.110 2.150 5.350 3.365 ;
        RECT  3.910 0.990 5.110 1.390 ;
        RECT  3.910 2.150 5.110 2.550 ;
        RECT  3.670 0.495 3.910 1.390 ;
        RECT  3.670 2.150 3.910 3.365 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 1.5138 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 1.800 2.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.480 -0.235 10.640 0.235 ;
        RECT  10.100 -0.235 10.480 1.215 ;
        RECT  9.040 -0.235 10.100 0.235 ;
        RECT  8.660 -0.235 9.040 0.745 ;
        RECT  7.580 -0.235 8.660 0.235 ;
        RECT  7.200 -0.235 7.580 0.745 ;
        RECT  6.140 -0.235 7.200 0.235 ;
        RECT  5.760 -0.235 6.140 0.745 ;
        RECT  4.700 -0.235 5.760 0.235 ;
        RECT  4.320 -0.235 4.700 0.745 ;
        RECT  3.250 -0.235 4.320 0.235 ;
        RECT  2.870 -0.235 3.250 1.255 ;
        RECT  1.820 -0.235 2.870 0.235 ;
        RECT  1.440 -0.235 1.820 0.740 ;
        RECT  0.475 -0.235 1.440 0.235 ;
        RECT  0.220 -0.235 0.475 0.535 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.480 3.685 10.640 4.155 ;
        RECT  10.100 2.300 10.480 4.155 ;
        RECT  9.040 3.685 10.100 4.155 ;
        RECT  8.660 2.780 9.040 4.155 ;
        RECT  7.580 3.685 8.660 4.155 ;
        RECT  7.200 2.780 7.580 4.155 ;
        RECT  6.140 3.685 7.200 4.155 ;
        RECT  5.760 2.780 6.140 4.155 ;
        RECT  4.700 3.685 5.760 4.155 ;
        RECT  4.320 2.780 4.700 4.155 ;
        RECT  3.250 3.685 4.320 4.155 ;
        RECT  2.870 2.305 3.250 4.155 ;
        RECT  1.820 3.685 2.870 4.155 ;
        RECT  1.440 2.935 1.820 4.155 ;
        RECT  0.475 3.685 1.440 4.155 ;
        RECT  0.230 3.390 0.475 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.450 0.495 9.690 1.390 ;
        RECT  9.450 2.150 9.690 3.365 ;
        RECT  8.230 0.990 9.450 1.390 ;
        RECT  8.230 2.150 9.450 2.550 ;
        RECT  7.990 0.495 8.230 1.390 ;
        RECT  7.990 2.150 8.230 3.365 ;
        RECT  7.650 0.990 7.990 1.390 ;
        RECT  7.650 2.150 7.990 2.550 ;
        RECT  5.350 0.990 5.790 1.390 ;
        RECT  5.350 2.150 5.790 2.550 ;
        RECT  5.110 0.495 5.350 1.390 ;
        RECT  5.110 2.150 5.350 3.365 ;
        RECT  3.910 0.990 5.110 1.390 ;
        RECT  3.910 2.150 5.110 2.550 ;
        RECT  3.670 0.495 3.910 1.390 ;
        RECT  3.670 2.150 3.910 3.365 ;
        RECT  2.470 1.620 5.195 1.920 ;
        RECT  2.230 0.495 2.470 3.380 ;
        RECT  0.740 1.010 2.230 1.255 ;
        RECT  0.730 2.440 2.230 2.670 ;
    END
END BUFFD10BWP7T

MACRO BUFFD12BWP7T
    CLASS CORE ;
    FOREIGN BUFFD12BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 7.7736 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.020 0.500 11.360 1.410 ;
        RECT  11.020 2.120 11.360 3.380 ;
        RECT  9.920 1.010 11.020 1.410 ;
        RECT  9.920 2.120 11.020 2.520 ;
        RECT  9.580 0.500 9.920 1.410 ;
        RECT  9.580 2.120 9.920 3.380 ;
        RECT  8.570 1.010 9.580 1.410 ;
        RECT  8.570 2.120 9.580 2.520 ;
        RECT  8.470 1.010 8.570 2.520 ;
        RECT  8.130 0.500 8.470 3.380 ;
        RECT  7.110 1.010 8.130 2.520 ;
        RECT  7.020 1.010 7.110 1.410 ;
        RECT  7.020 2.120 7.110 2.520 ;
        RECT  6.680 0.500 7.020 1.410 ;
        RECT  6.680 2.120 7.020 3.380 ;
        RECT  5.560 1.010 6.680 1.410 ;
        RECT  5.560 2.120 6.680 2.520 ;
        RECT  5.220 0.500 5.560 1.410 ;
        RECT  5.220 2.120 5.560 3.380 ;
        RECT  4.120 1.010 5.220 1.410 ;
        RECT  4.120 2.120 5.220 2.520 ;
        RECT  3.780 0.500 4.120 1.410 ;
        RECT  3.780 2.120 4.120 3.380 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.650 1.605 2.040 2.100 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.120 -0.235 12.320 0.235 ;
        RECT  11.780 -0.235 12.120 1.195 ;
        RECT  10.640 -0.235 11.780 0.235 ;
        RECT  10.300 -0.235 10.640 0.760 ;
        RECT  9.190 -0.235 10.300 0.235 ;
        RECT  8.850 -0.235 9.190 0.760 ;
        RECT  7.740 -0.235 8.850 0.235 ;
        RECT  7.400 -0.235 7.740 0.760 ;
        RECT  6.280 -0.235 7.400 0.235 ;
        RECT  5.940 -0.235 6.280 0.760 ;
        RECT  4.840 -0.235 5.940 0.235 ;
        RECT  4.500 -0.235 4.840 0.760 ;
        RECT  3.400 -0.235 4.500 0.235 ;
        RECT  3.060 -0.235 3.400 1.200 ;
        RECT  1.960 -0.235 3.060 0.235 ;
        RECT  1.620 -0.235 1.960 0.760 ;
        RECT  0.520 -0.235 1.620 0.235 ;
        RECT  0.180 -0.235 0.520 1.200 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.120 3.685 12.320 4.155 ;
        RECT  11.780 2.305 12.120 4.155 ;
        RECT  10.640 3.685 11.780 4.155 ;
        RECT  10.300 2.750 10.640 4.155 ;
        RECT  9.190 3.685 10.300 4.155 ;
        RECT  8.850 2.750 9.190 4.155 ;
        RECT  7.740 3.685 8.850 4.155 ;
        RECT  7.400 2.750 7.740 4.155 ;
        RECT  6.280 3.685 7.400 4.155 ;
        RECT  5.940 2.750 6.280 4.155 ;
        RECT  4.840 3.685 5.940 4.155 ;
        RECT  4.500 2.750 4.840 4.155 ;
        RECT  3.400 3.685 4.500 4.155 ;
        RECT  3.060 2.310 3.400 4.155 ;
        RECT  1.960 3.685 3.060 4.155 ;
        RECT  1.620 2.850 1.960 4.155 ;
        RECT  0.470 3.685 1.620 4.155 ;
        RECT  0.230 2.480 0.470 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.020 0.500 11.360 1.410 ;
        RECT  11.020 2.120 11.360 3.380 ;
        RECT  9.920 1.010 11.020 1.410 ;
        RECT  9.920 2.120 11.020 2.520 ;
        RECT  9.580 0.500 9.920 1.410 ;
        RECT  9.580 2.120 9.920 3.380 ;
        RECT  8.770 1.010 9.580 1.410 ;
        RECT  8.770 2.120 9.580 2.520 ;
        RECT  6.680 0.500 6.910 1.410 ;
        RECT  6.680 2.120 6.910 3.380 ;
        RECT  5.560 1.010 6.680 1.410 ;
        RECT  5.560 2.120 6.680 2.520 ;
        RECT  5.220 0.500 5.560 1.410 ;
        RECT  5.220 2.120 5.560 3.380 ;
        RECT  4.120 1.010 5.220 1.410 ;
        RECT  4.120 2.120 5.220 2.520 ;
        RECT  3.780 0.500 4.120 1.410 ;
        RECT  3.780 2.120 4.120 3.380 ;
        RECT  2.680 1.640 6.820 1.890 ;
        RECT  2.340 0.500 2.680 3.380 ;
        RECT  1.240 1.025 2.340 1.255 ;
        RECT  1.240 2.380 2.340 2.610 ;
        RECT  0.900 0.500 1.240 1.255 ;
        RECT  0.900 2.380 1.240 3.380 ;
    END
END BUFFD12BWP7T

MACRO BUFFD1BWP7T
    CLASS CORE ;
    FOREIGN BUFFD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1731 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.775 0.495 2.100 3.415 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.660 0.980 2.710 ;
        RECT  0.630 1.660 0.700 2.000 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.350 -0.235 2.240 0.235 ;
        RECT  0.970 -0.235 1.350 0.880 ;
        RECT  0.000 -0.235 0.970 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.350 3.685 2.240 4.155 ;
        RECT  0.970 2.990 1.350 4.155 ;
        RECT  0.000 3.685 0.970 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.315 1.120 1.545 2.000 ;
        RECT  0.470 1.120 1.315 1.380 ;
        RECT  0.400 0.965 0.470 1.380 ;
        RECT  0.400 2.335 0.470 2.685 ;
        RECT  0.170 0.965 0.400 2.685 ;
    END
END BUFFD1BWP7T

MACRO BUFFD1P5BWP7T
    CLASS CORE ;
    FOREIGN BUFFD1P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.0114 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.995 2.660 2.720 ;
        RECT  1.585 0.995 2.380 1.230 ;
        RECT  1.675 2.370 2.380 2.720 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.640 1.210 0.980 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 -0.235 2.800 0.235 ;
        RECT  2.325 -0.235 2.570 0.535 ;
        RECT  1.260 -0.235 2.325 0.235 ;
        RECT  0.900 -0.235 1.260 0.935 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 3.685 2.800 4.155 ;
        RECT  2.320 3.230 2.575 4.155 ;
        RECT  1.250 3.685 2.320 4.155 ;
        RECT  0.885 3.075 1.250 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.445 1.605 2.135 1.955 ;
        RECT  1.215 1.605 1.445 2.835 ;
        RECT  0.470 2.595 1.215 2.835 ;
        RECT  0.370 0.515 0.525 0.755 ;
        RECT  0.370 2.595 0.470 3.370 ;
        RECT  0.230 0.515 0.370 3.370 ;
        RECT  0.140 0.515 0.230 2.835 ;
    END
END BUFFD1P5BWP7T

MACRO BUFFD2BWP7T
    CLASS CORE ;
    FOREIGN BUFFD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.5642 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.090 2.660 2.580 ;
        RECT  2.170 1.090 2.380 1.370 ;
        RECT  2.160 2.340 2.380 2.580 ;
        RECT  1.930 0.495 2.170 1.370 ;
        RECT  1.925 2.340 2.160 3.390 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.480 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.235 3.360 0.235 ;
        RECT  2.890 -0.235 3.125 1.255 ;
        RECT  1.440 -0.235 2.890 0.235 ;
        RECT  1.190 -0.235 1.440 1.255 ;
        RECT  0.000 -0.235 1.190 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 3.685 3.360 4.155 ;
        RECT  2.895 2.250 3.125 4.155 ;
        RECT  1.430 3.685 2.895 4.155 ;
        RECT  1.190 2.250 1.430 4.155 ;
        RECT  0.000 3.685 1.190 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.960 1.660 2.150 1.895 ;
        RECT  0.720 1.070 0.960 3.240 ;
        RECT  0.530 1.070 0.720 1.310 ;
        RECT  0.240 3.000 0.720 3.240 ;
        RECT  0.290 0.495 0.530 1.310 ;
    END
END BUFFD2BWP7T

MACRO BUFFD2P5BWP7T
    CLASS CORE ;
    FOREIGN BUFFD2P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.1093 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 0.515 3.740 1.335 ;
        RECT  3.530 2.205 3.685 3.395 ;
        RECT  3.455 0.515 3.530 3.395 ;
        RECT  3.400 0.515 3.455 2.555 ;
        RECT  2.640 0.985 3.400 2.555 ;
        RECT  2.190 0.985 2.640 1.335 ;
        RECT  2.195 2.205 2.640 2.555 ;
        RECT  1.960 2.205 2.195 3.375 ;
        RECT  1.950 0.495 2.190 1.335 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.480 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 -0.235 3.920 0.235 ;
        RECT  2.660 -0.235 3.040 0.735 ;
        RECT  1.420 -0.235 2.660 0.235 ;
        RECT  1.170 -0.235 1.420 1.255 ;
        RECT  0.000 -0.235 1.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 3.685 3.920 4.155 ;
        RECT  2.660 2.985 3.040 4.155 ;
        RECT  1.410 3.685 2.660 4.155 ;
        RECT  1.170 2.250 1.410 4.155 ;
        RECT  0.000 3.685 1.170 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.940 1.660 2.350 1.895 ;
        RECT  0.710 1.070 0.940 3.240 ;
        RECT  0.530 1.070 0.710 1.310 ;
        RECT  0.240 3.000 0.710 3.240 ;
        RECT  0.290 0.495 0.530 1.310 ;
    END
END BUFFD2P5BWP7T

MACRO BUFFD3BWP7T
    CLASS CORE ;
    FOREIGN BUFFD3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.6781 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 0.475 3.685 1.335 ;
        RECT  3.530 2.155 3.685 3.385 ;
        RECT  3.455 0.475 3.530 3.385 ;
        RECT  2.640 0.985 3.455 2.505 ;
        RECT  2.190 0.985 2.640 1.335 ;
        RECT  2.195 2.155 2.640 2.505 ;
        RECT  1.960 2.155 2.195 3.385 ;
        RECT  1.950 0.495 2.190 1.335 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.480 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 -0.235 3.920 0.235 ;
        RECT  2.660 -0.235 3.040 0.735 ;
        RECT  1.420 -0.235 2.660 0.235 ;
        RECT  1.170 -0.235 1.420 1.255 ;
        RECT  0.000 -0.235 1.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 3.685 3.920 4.155 ;
        RECT  2.660 2.780 3.040 4.155 ;
        RECT  1.410 3.685 2.660 4.155 ;
        RECT  1.170 2.250 1.410 4.155 ;
        RECT  0.000 3.685 1.170 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.940 1.660 2.370 1.895 ;
        RECT  0.710 1.070 0.940 3.240 ;
        RECT  0.530 1.070 0.710 1.310 ;
        RECT  0.240 3.000 0.710 3.240 ;
        RECT  0.290 0.495 0.530 1.310 ;
    END
END BUFFD3BWP7T

MACRO BUFFD4BWP7T
    CLASS CORE ;
    FOREIGN BUFFD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.855 0.475 4.090 3.430 ;
        RECT  3.190 0.985 3.855 2.505 ;
        RECT  2.650 0.985 3.190 1.335 ;
        RECT  2.650 2.155 3.190 2.505 ;
        RECT  2.410 0.495 2.650 1.335 ;
        RECT  2.415 2.155 2.650 3.430 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.480 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 -0.235 5.040 0.235 ;
        RECT  4.500 -0.235 4.880 1.205 ;
        RECT  3.440 -0.235 4.500 0.235 ;
        RECT  3.060 -0.235 3.440 0.735 ;
        RECT  1.990 -0.235 3.060 0.235 ;
        RECT  1.610 -0.235 1.990 1.205 ;
        RECT  0.540 -0.235 1.610 0.235 ;
        RECT  0.160 -0.235 0.540 1.205 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 3.685 5.040 4.155 ;
        RECT  4.500 2.305 4.880 4.155 ;
        RECT  3.440 3.685 4.500 4.155 ;
        RECT  3.060 2.780 3.440 4.155 ;
        RECT  1.990 3.685 3.060 4.155 ;
        RECT  1.610 2.305 1.990 4.155 ;
        RECT  0.540 3.685 1.610 4.155 ;
        RECT  0.160 2.940 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.650 0.985 2.990 1.335 ;
        RECT  2.650 2.155 2.990 2.505 ;
        RECT  2.410 0.495 2.650 1.335 ;
        RECT  2.415 2.155 2.650 3.430 ;
        RECT  1.185 1.660 2.930 1.895 ;
        RECT  0.955 0.495 1.185 3.430 ;
    END
END BUFFD4BWP7T

MACRO BUFFD5BWP7T
    CLASS CORE ;
    FOREIGN BUFFD5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 3.8157 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.475 0.470 5.710 1.335 ;
        RECT  5.475 2.155 5.710 3.405 ;
        RECT  4.650 0.985 5.475 1.335 ;
        RECT  4.650 2.155 5.475 2.505 ;
        RECT  4.210 0.985 4.650 2.505 ;
        RECT  3.975 0.470 4.210 3.405 ;
        RECT  3.750 0.985 3.975 2.505 ;
        RECT  2.710 0.985 3.750 1.335 ;
        RECT  2.710 2.155 3.750 2.505 ;
        RECT  2.470 0.490 2.710 1.335 ;
        RECT  2.475 2.155 2.710 3.405 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.480 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.030 -0.235 6.160 0.235 ;
        RECT  4.650 -0.235 5.030 0.735 ;
        RECT  3.530 -0.235 4.650 0.235 ;
        RECT  3.150 -0.235 3.530 0.735 ;
        RECT  2.030 -0.235 3.150 0.235 ;
        RECT  1.650 -0.235 2.030 1.205 ;
        RECT  0.560 -0.235 1.650 0.235 ;
        RECT  0.180 -0.235 0.560 1.205 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.030 3.685 6.160 4.155 ;
        RECT  4.650 2.780 5.030 4.155 ;
        RECT  3.530 3.685 4.650 4.155 ;
        RECT  3.150 2.780 3.530 4.155 ;
        RECT  2.030 3.685 3.150 4.155 ;
        RECT  1.650 2.305 2.030 4.155 ;
        RECT  0.560 3.685 1.650 4.155 ;
        RECT  0.180 2.940 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.475 0.470 5.710 1.335 ;
        RECT  5.475 2.155 5.710 3.405 ;
        RECT  4.850 0.985 5.475 1.335 ;
        RECT  4.850 2.155 5.475 2.505 ;
        RECT  2.710 0.985 3.550 1.335 ;
        RECT  2.710 2.155 3.550 2.505 ;
        RECT  2.470 0.490 2.710 1.335 ;
        RECT  2.475 2.155 2.710 3.405 ;
        RECT  1.205 1.660 3.460 1.895 ;
        RECT  0.975 0.495 1.205 3.405 ;
    END
END BUFFD5BWP7T

MACRO BUFFD6BWP7T
    CLASS CORE ;
    FOREIGN BUFFD6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 3.8394 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.295 0.475 5.530 1.335 ;
        RECT  5.295 2.155 5.530 3.420 ;
        RECT  4.650 0.985 5.295 1.335 ;
        RECT  4.650 2.155 5.295 2.505 ;
        RECT  4.090 0.985 4.650 2.505 ;
        RECT  3.855 0.475 4.090 3.420 ;
        RECT  3.750 0.985 3.855 2.505 ;
        RECT  2.650 0.985 3.750 1.335 ;
        RECT  2.650 2.155 3.750 2.505 ;
        RECT  2.410 0.495 2.650 1.335 ;
        RECT  2.415 2.155 2.650 3.420 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.480 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.340 -0.235 6.720 0.235 ;
        RECT  5.960 -0.235 6.340 1.205 ;
        RECT  4.880 -0.235 5.960 0.235 ;
        RECT  4.500 -0.235 4.880 0.735 ;
        RECT  3.440 -0.235 4.500 0.235 ;
        RECT  3.060 -0.235 3.440 0.735 ;
        RECT  1.990 -0.235 3.060 0.235 ;
        RECT  1.610 -0.235 1.990 1.205 ;
        RECT  0.540 -0.235 1.610 0.235 ;
        RECT  0.160 -0.235 0.540 1.205 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.340 3.685 6.720 4.155 ;
        RECT  5.960 2.305 6.340 4.155 ;
        RECT  4.880 3.685 5.960 4.155 ;
        RECT  4.500 2.780 4.880 4.155 ;
        RECT  3.440 3.685 4.500 4.155 ;
        RECT  3.060 2.780 3.440 4.155 ;
        RECT  1.990 3.685 3.060 4.155 ;
        RECT  1.610 2.305 1.990 4.155 ;
        RECT  0.540 3.685 1.610 4.155 ;
        RECT  0.160 2.950 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.295 0.475 5.530 1.335 ;
        RECT  5.295 2.155 5.530 3.420 ;
        RECT  4.850 0.985 5.295 1.335 ;
        RECT  4.850 2.155 5.295 2.505 ;
        RECT  2.650 0.985 3.550 1.335 ;
        RECT  2.650 2.155 3.550 2.505 ;
        RECT  2.410 0.495 2.650 1.335 ;
        RECT  2.415 2.155 2.650 3.420 ;
        RECT  1.185 1.660 3.400 1.895 ;
        RECT  0.955 0.495 1.185 3.420 ;
    END
END BUFFD6BWP7T

MACRO BUFFD8BWP7T
    CLASS CORE ;
    FOREIGN BUFFD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 5.1192 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.430 0.495 7.670 1.365 ;
        RECT  7.430 2.150 7.665 3.435 ;
        RECT  6.330 1.015 7.430 1.365 ;
        RECT  6.330 2.150 7.430 2.550 ;
        RECT  6.225 1.015 6.330 2.550 ;
        RECT  5.990 0.475 6.225 3.435 ;
        RECT  5.430 1.015 5.990 2.550 ;
        RECT  4.790 1.015 5.430 1.365 ;
        RECT  4.790 2.150 5.430 2.550 ;
        RECT  4.555 0.475 4.790 1.365 ;
        RECT  4.555 2.150 4.790 3.435 ;
        RECT  3.350 1.015 4.555 1.365 ;
        RECT  3.350 2.150 4.555 2.550 ;
        RECT  3.110 0.495 3.350 1.365 ;
        RECT  3.115 2.150 3.350 3.435 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.650 1.400 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.460 -0.235 8.960 0.235 ;
        RECT  8.080 -0.235 8.460 1.205 ;
        RECT  7.020 -0.235 8.080 0.235 ;
        RECT  6.640 -0.235 7.020 0.735 ;
        RECT  5.580 -0.235 6.640 0.235 ;
        RECT  5.200 -0.235 5.580 0.735 ;
        RECT  4.140 -0.235 5.200 0.235 ;
        RECT  3.760 -0.235 4.140 0.735 ;
        RECT  2.700 -0.235 3.760 0.235 ;
        RECT  2.320 -0.235 2.700 1.205 ;
        RECT  1.260 -0.235 2.320 0.235 ;
        RECT  0.880 -0.235 1.260 0.785 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.460 3.685 8.960 4.155 ;
        RECT  8.080 2.305 8.460 4.155 ;
        RECT  7.020 3.685 8.080 4.155 ;
        RECT  6.640 2.780 7.020 4.155 ;
        RECT  5.580 3.685 6.640 4.155 ;
        RECT  5.200 2.780 5.580 4.155 ;
        RECT  4.140 3.685 5.200 4.155 ;
        RECT  3.760 2.780 4.140 4.155 ;
        RECT  2.700 3.685 3.760 4.155 ;
        RECT  2.320 2.305 2.700 4.155 ;
        RECT  1.260 3.685 2.320 4.155 ;
        RECT  0.880 2.980 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.430 0.495 7.670 1.365 ;
        RECT  7.430 2.150 7.665 3.435 ;
        RECT  6.530 1.015 7.430 1.365 ;
        RECT  6.530 2.150 7.430 2.550 ;
        RECT  4.790 1.015 5.230 1.365 ;
        RECT  4.790 2.150 5.230 2.550 ;
        RECT  4.555 0.475 4.790 1.365 ;
        RECT  4.555 2.150 4.790 3.435 ;
        RECT  3.350 1.015 4.555 1.365 ;
        RECT  3.350 2.150 4.555 2.550 ;
        RECT  3.110 0.495 3.350 1.365 ;
        RECT  3.115 2.150 3.350 3.435 ;
        RECT  1.905 1.615 5.040 1.920 ;
        RECT  1.675 0.495 1.905 3.435 ;
        RECT  0.465 1.075 1.675 1.305 ;
        RECT  0.470 2.510 1.675 2.740 ;
        RECT  0.230 2.510 0.470 3.320 ;
        RECT  0.235 0.495 0.465 1.305 ;
    END
END BUFFD8BWP7T

MACRO BUFTD0BWP7T
    CLASS CORE ;
    FOREIGN BUFTD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5560 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.420 5.460 3.285 ;
        RECT  4.650 1.420 5.180 1.660 ;
        RECT  5.055 3.040 5.180 3.285 ;
        RECT  4.410 0.965 4.650 1.660 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 1.500 3.620 2.670 ;
        RECT  2.990 2.430 3.380 2.670 ;
        RECT  2.750 2.430 2.990 3.210 ;
        RECT  0.980 2.980 2.750 3.210 ;
        RECT  0.700 1.770 0.980 3.210 ;
        RECT  0.630 1.770 0.700 2.160 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.590 2.935 1.830 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.125 1.590 2.380 1.830 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.440 -0.235 5.600 0.235 ;
        RECT  5.060 -0.235 5.440 1.170 ;
        RECT  2.720 -0.235 5.060 0.235 ;
        RECT  2.380 -0.235 2.720 0.470 ;
        RECT  1.260 -0.235 2.380 0.235 ;
        RECT  0.880 -0.235 1.260 0.825 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.590 3.685 5.600 4.155 ;
        RECT  4.350 2.990 4.590 4.155 ;
        RECT  2.860 3.685 4.350 4.155 ;
        RECT  2.520 3.450 2.860 4.155 ;
        RECT  1.080 3.685 2.520 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.110 2.080 4.910 2.320 ;
        RECT  3.325 0.465 4.345 0.695 ;
        RECT  3.870 1.020 4.110 3.280 ;
        RECT  3.660 1.020 3.870 1.250 ;
        RECT  3.420 3.040 3.870 3.280 ;
        RECT  3.085 0.465 3.325 0.980 ;
        RECT  1.910 0.740 3.085 0.980 ;
        RECT  1.895 2.490 2.450 2.730 ;
        RECT  1.895 0.540 1.910 0.980 ;
        RECT  1.655 0.540 1.895 2.730 ;
        RECT  0.465 1.120 1.380 1.460 ;
        RECT  0.370 0.560 0.465 1.460 ;
        RECT  0.370 2.495 0.465 2.835 ;
        RECT  0.140 0.560 0.370 2.835 ;
    END
END BUFTD0BWP7T

MACRO BUFTD1BWP7T
    CLASS CORE ;
    FOREIGN BUFTD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.9488 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 1.220 5.460 2.830 ;
        RECT  5.180 1.220 5.345 3.290 ;
        RECT  4.650 1.220 5.180 1.460 ;
        RECT  5.105 2.245 5.180 3.290 ;
        RECT  4.410 0.965 4.650 1.460 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.4626 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 1.500 3.620 2.670 ;
        RECT  2.990 2.430 3.380 2.670 ;
        RECT  2.750 2.430 2.990 3.210 ;
        RECT  0.980 2.980 2.750 3.210 ;
        RECT  0.700 1.770 0.980 3.210 ;
        RECT  0.630 1.770 0.700 2.160 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.5760 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.590 2.935 1.830 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.125 1.590 2.380 1.830 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.440 -0.235 5.600 0.235 ;
        RECT  5.060 -0.235 5.440 0.980 ;
        RECT  2.720 -0.235 5.060 0.235 ;
        RECT  2.380 -0.235 2.720 0.470 ;
        RECT  1.260 -0.235 2.380 0.235 ;
        RECT  0.880 -0.235 1.260 0.825 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.590 3.685 5.600 4.155 ;
        RECT  4.350 2.245 4.590 4.155 ;
        RECT  3.000 3.685 4.350 4.155 ;
        RECT  2.660 3.450 3.000 4.155 ;
        RECT  1.080 3.685 2.660 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.110 1.755 4.420 1.995 ;
        RECT  3.325 0.465 4.340 0.695 ;
        RECT  3.870 1.020 4.110 3.345 ;
        RECT  3.660 1.020 3.870 1.250 ;
        RECT  3.420 3.105 3.870 3.345 ;
        RECT  3.085 0.465 3.325 0.980 ;
        RECT  1.910 0.750 3.085 0.980 ;
        RECT  1.895 2.490 2.450 2.730 ;
        RECT  1.895 0.540 1.910 0.980 ;
        RECT  1.655 0.540 1.895 2.730 ;
        RECT  0.465 1.120 1.380 1.460 ;
        RECT  0.370 0.540 0.465 1.460 ;
        RECT  0.370 2.425 0.465 2.765 ;
        RECT  0.140 0.540 0.370 2.765 ;
    END
END BUFTD1BWP7T

MACRO BUFTD2BWP7T
    CLASS CORE ;
    FOREIGN BUFTD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.0800 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.020 6.020 2.740 ;
        RECT  5.205 1.020 5.740 1.260 ;
        RECT  5.185 2.440 5.740 2.740 ;
        RECT  4.975 0.620 5.205 1.260 ;
        RECT  4.945 2.440 5.185 3.410 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.4536 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.385 1.760 3.625 2.670 ;
        RECT  2.965 2.430 3.385 2.670 ;
        RECT  2.725 2.430 2.965 3.220 ;
        RECT  0.980 2.980 2.725 3.220 ;
        RECT  0.700 1.770 0.980 3.220 ;
        RECT  0.610 1.770 0.700 2.120 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.5517 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.675 2.955 1.915 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.145 1.675 2.380 1.915 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.000 -0.235 6.160 0.235 ;
        RECT  5.620 -0.235 6.000 0.785 ;
        RECT  4.500 -0.235 5.620 0.235 ;
        RECT  4.160 -0.235 4.500 0.470 ;
        RECT  2.735 -0.235 4.160 0.235 ;
        RECT  2.315 -0.235 2.735 0.465 ;
        RECT  1.260 -0.235 2.315 0.235 ;
        RECT  0.880 -0.235 1.260 0.825 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.000 3.685 6.160 4.155 ;
        RECT  5.620 3.050 6.000 4.155 ;
        RECT  4.475 3.685 5.620 4.155 ;
        RECT  4.135 3.455 4.475 4.155 ;
        RECT  2.895 3.685 4.135 4.155 ;
        RECT  2.555 3.450 2.895 4.155 ;
        RECT  1.060 3.685 2.555 4.155 ;
        RECT  0.720 3.455 1.060 4.155 ;
        RECT  0.000 3.685 0.720 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.745 1.510 5.455 1.750 ;
        RECT  4.505 0.700 4.745 1.750 ;
        RECT  1.905 0.700 4.505 0.930 ;
        RECT  4.105 1.890 4.290 2.230 ;
        RECT  3.875 1.160 4.105 3.225 ;
        RECT  3.595 1.160 3.875 1.390 ;
        RECT  3.375 2.985 3.875 3.225 ;
        RECT  1.905 2.510 2.355 2.750 ;
        RECT  1.675 0.580 1.905 2.750 ;
        RECT  0.465 1.120 1.375 1.460 ;
        RECT  0.380 2.440 0.470 2.780 ;
        RECT  0.380 0.540 0.465 1.460 ;
        RECT  0.140 0.540 0.380 2.780 ;
    END
END BUFTD2BWP7T

MACRO BUFTD3BWP7T
    CLASS CORE ;
    FOREIGN BUFTD3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.1467 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  6.890 0.580 7.055 1.285 ;
        RECT  6.890 2.380 7.050 3.410 ;
        RECT  6.810 0.580 6.890 3.410 ;
        RECT  5.990 1.015 6.810 2.730 ;
        RECT  5.610 1.015 5.990 1.285 ;
        RECT  5.525 2.380 5.990 2.730 ;
        RECT  5.370 0.700 5.610 1.285 ;
        RECT  5.285 2.380 5.525 3.410 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.4599 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 1.620 3.645 2.670 ;
        RECT  2.965 2.430 3.405 2.670 ;
        RECT  2.725 2.430 2.965 3.220 ;
        RECT  0.980 2.980 2.725 3.220 ;
        RECT  0.700 1.770 0.980 3.220 ;
        RECT  0.610 1.770 0.700 2.120 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.5580 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.720 2.955 1.960 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.145 1.720 2.380 1.960 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.400 -0.235 7.280 0.235 ;
        RECT  6.020 -0.235 6.400 0.785 ;
        RECT  4.850 -0.235 6.020 0.235 ;
        RECT  4.485 -0.235 4.850 0.465 ;
        RECT  2.720 -0.235 4.485 0.235 ;
        RECT  2.380 -0.235 2.720 0.465 ;
        RECT  1.260 -0.235 2.380 0.235 ;
        RECT  0.880 -0.235 1.260 0.825 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.375 3.685 7.280 4.155 ;
        RECT  5.995 2.980 6.375 4.155 ;
        RECT  4.705 3.685 5.995 4.155 ;
        RECT  4.365 2.555 4.705 4.155 ;
        RECT  3.075 3.685 4.365 4.155 ;
        RECT  2.735 3.450 3.075 4.155 ;
        RECT  1.060 3.685 2.735 4.155 ;
        RECT  0.720 3.455 1.060 4.155 ;
        RECT  0.000 3.685 0.720 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.610 1.015 5.790 1.285 ;
        RECT  5.525 2.380 5.790 2.730 ;
        RECT  5.370 0.700 5.610 1.285 ;
        RECT  5.065 1.515 5.455 1.750 ;
        RECT  4.825 0.695 5.065 1.750 ;
        RECT  1.905 0.695 4.825 0.925 ;
        RECT  4.120 1.945 4.630 2.180 ;
        RECT  3.890 1.155 4.120 3.350 ;
        RECT  3.780 1.155 3.890 1.385 ;
        RECT  3.495 3.120 3.890 3.350 ;
        RECT  1.905 2.510 2.375 2.750 ;
        RECT  1.675 0.580 1.905 2.750 ;
        RECT  0.465 1.120 1.375 1.460 ;
        RECT  0.380 2.440 0.470 2.780 ;
        RECT  0.380 0.540 0.465 1.460 ;
        RECT  0.140 0.540 0.380 2.780 ;
        RECT  5.285 2.380 5.525 3.410 ;
    END
END BUFTD3BWP7T

MACRO BUFTD4BWP7T
    CLASS CORE ;
    FOREIGN BUFTD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.1708 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  6.640 0.615 6.890 3.410 ;
        RECT  6.610 1.020 6.640 3.410 ;
        RECT  5.990 1.020 6.610 2.740 ;
        RECT  5.440 1.020 5.990 1.260 ;
        RECT  5.410 2.440 5.990 2.740 ;
        RECT  5.195 0.615 5.440 1.260 ;
        RECT  5.170 2.440 5.410 3.410 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.4599 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 1.620 3.645 2.670 ;
        RECT  2.965 2.430 3.405 2.670 ;
        RECT  2.725 2.430 2.965 3.220 ;
        RECT  0.980 2.980 2.725 3.220 ;
        RECT  0.700 1.770 0.980 3.220 ;
        RECT  0.610 1.770 0.700 2.120 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 0.5580 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.720 2.955 1.960 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.145 1.720 2.380 1.960 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.665 -0.235 7.840 0.235 ;
        RECT  7.285 -0.235 7.665 0.905 ;
        RECT  6.225 -0.235 7.285 0.235 ;
        RECT  5.845 -0.235 6.225 0.785 ;
        RECT  4.695 -0.235 5.845 0.235 ;
        RECT  4.275 -0.235 4.695 0.465 ;
        RECT  2.720 -0.235 4.275 0.235 ;
        RECT  2.380 -0.235 2.720 0.465 ;
        RECT  1.260 -0.235 2.380 0.235 ;
        RECT  0.880 -0.235 1.260 0.825 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.640 3.685 7.840 4.155 ;
        RECT  7.260 2.590 7.640 4.155 ;
        RECT  6.200 3.685 7.260 4.155 ;
        RECT  5.820 3.000 6.200 4.155 ;
        RECT  4.750 3.685 5.820 4.155 ;
        RECT  4.370 2.555 4.750 4.155 ;
        RECT  3.075 3.685 4.370 4.155 ;
        RECT  2.735 3.450 3.075 4.155 ;
        RECT  1.060 3.685 2.735 4.155 ;
        RECT  0.720 3.455 1.060 4.155 ;
        RECT  0.000 3.685 0.720 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.440 1.020 5.790 1.260 ;
        RECT  5.410 2.440 5.790 2.740 ;
        RECT  5.195 0.615 5.440 1.260 ;
        RECT  5.170 2.440 5.410 3.410 ;
        RECT  4.725 0.695 4.965 1.750 ;
        RECT  1.905 0.695 4.725 0.925 ;
        RECT  4.120 1.890 4.495 2.230 ;
        RECT  3.890 1.155 4.120 3.350 ;
        RECT  3.595 1.155 3.890 1.385 ;
        RECT  3.495 3.120 3.890 3.350 ;
        RECT  1.905 2.510 2.375 2.750 ;
        RECT  1.675 0.580 1.905 2.750 ;
        RECT  0.465 1.120 1.375 1.460 ;
        RECT  0.380 2.440 0.470 2.780 ;
        RECT  0.380 0.540 0.465 1.460 ;
        RECT  0.140 0.540 0.380 2.780 ;
        RECT  4.965 1.510 5.680 1.750 ;
    END
END BUFTD4BWP7T

MACRO BUFTD6BWP7T
    CLASS CORE ;
    FOREIGN BUFTD6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 3.4020 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  10.000 0.635 10.250 1.300 ;
        RECT  10.005 2.380 10.245 3.380 ;
        RECT  9.690 2.380 10.005 2.730 ;
        RECT  9.690 1.020 10.000 1.300 ;
        RECT  8.805 1.020 9.690 2.730 ;
        RECT  8.790 0.635 8.805 3.380 ;
        RECT  8.565 0.635 8.790 1.300 ;
        RECT  8.565 2.380 8.790 3.380 ;
        RECT  7.365 1.020 8.565 1.300 ;
        RECT  7.365 2.380 8.565 2.730 ;
        RECT  7.125 0.680 7.365 1.300 ;
        RECT  7.125 2.380 7.365 3.380 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.7353 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.760 2.020 4.990 2.755 ;
        RECT  3.885 2.515 4.760 2.755 ;
        RECT  3.645 2.515 3.885 3.225 ;
        RECT  3.090 2.985 3.645 3.225 ;
        RECT  2.860 2.985 3.090 3.455 ;
        RECT  1.760 3.225 2.860 3.455 ;
        RECT  1.530 2.940 1.760 3.455 ;
        RECT  1.030 2.940 1.530 3.170 ;
        RECT  0.980 2.650 1.030 3.170 ;
        RECT  0.800 1.615 0.980 3.170 ;
        RECT  0.650 1.615 0.800 3.030 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 1.1574 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 1.595 3.860 1.825 ;
        RECT  2.715 1.595 2.945 2.285 ;
        RECT  1.720 2.055 2.715 2.285 ;
        RECT  1.540 1.585 1.720 2.285 ;
        RECT  1.260 1.585 1.540 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 -0.235 11.200 0.235 ;
        RECT  10.655 -0.235 11.035 0.930 ;
        RECT  9.590 -0.235 10.655 0.235 ;
        RECT  9.210 -0.235 9.590 0.790 ;
        RECT  8.150 -0.235 9.210 0.235 ;
        RECT  7.770 -0.235 8.150 0.790 ;
        RECT  6.670 -0.235 7.770 0.235 ;
        RECT  6.330 -0.235 6.670 0.715 ;
        RECT  3.420 -0.235 6.330 0.235 ;
        RECT  3.040 -0.235 3.420 0.465 ;
        RECT  1.260 -0.235 3.040 0.235 ;
        RECT  0.880 -0.235 1.260 0.710 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.685 11.200 4.155 ;
        RECT  10.655 2.570 11.035 4.155 ;
        RECT  9.595 3.685 10.655 4.155 ;
        RECT  9.215 3.030 9.595 4.155 ;
        RECT  8.155 3.685 9.215 4.155 ;
        RECT  7.775 3.030 8.155 4.155 ;
        RECT  6.695 3.685 7.775 4.155 ;
        RECT  6.315 3.005 6.695 4.155 ;
        RECT  5.180 3.685 6.315 4.155 ;
        RECT  4.840 3.455 5.180 4.155 ;
        RECT  3.660 3.685 4.840 4.155 ;
        RECT  3.320 3.455 3.660 4.155 ;
        RECT  1.280 3.685 3.320 4.155 ;
        RECT  0.940 3.440 1.280 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.000 0.635 10.250 1.300 ;
        RECT  10.005 2.380 10.245 3.380 ;
        RECT  9.890 2.380 10.005 2.730 ;
        RECT  9.890 1.020 10.000 1.300 ;
        RECT  8.565 0.635 8.590 1.300 ;
        RECT  8.565 2.380 8.590 3.380 ;
        RECT  7.365 1.020 8.565 1.300 ;
        RECT  7.365 2.380 8.565 2.730 ;
        RECT  7.125 0.680 7.365 1.300 ;
        RECT  7.125 2.380 7.365 3.380 ;
        RECT  7.615 1.880 7.955 2.140 ;
        RECT  5.890 1.910 7.615 2.140 ;
        RECT  6.080 1.430 6.935 1.665 ;
        RECT  5.850 0.465 6.080 1.665 ;
        RECT  5.650 1.910 5.890 3.455 ;
        RECT  4.380 0.465 5.850 0.695 ;
        RECT  5.605 1.910 5.650 2.140 ;
        RECT  4.365 2.985 5.650 3.225 ;
        RECT  5.365 1.020 5.605 2.140 ;
        RECT  5.005 1.020 5.365 1.250 ;
        RECT  4.150 0.465 4.380 2.285 ;
        RECT  4.135 2.985 4.365 3.455 ;
        RECT  4.140 0.935 4.150 2.285 ;
        RECT  2.810 0.935 4.140 1.165 ;
        RECT  3.415 2.055 4.140 2.285 ;
        RECT  3.175 2.055 3.415 2.755 ;
        RECT  2.630 2.515 3.175 2.755 ;
        RECT  2.580 0.465 2.810 1.165 ;
        RECT  2.400 2.515 2.630 2.995 ;
        RECT  1.620 0.465 2.580 0.695 ;
        RECT  2.350 1.485 2.485 1.825 ;
        RECT  2.130 2.765 2.400 2.995 ;
        RECT  2.120 1.105 2.350 1.825 ;
        RECT  0.465 1.105 2.120 1.335 ;
        RECT  0.350 3.225 0.520 3.455 ;
        RECT  0.350 0.465 0.465 1.335 ;
        RECT  0.120 0.465 0.350 3.455 ;
    END
END BUFTD6BWP7T

MACRO BUFTD8BWP7T
    CLASS CORE ;
    FOREIGN BUFTD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 4.5360 ;
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  11.685 0.690 11.935 1.420 ;
        RECT  11.690 2.380 11.930 3.380 ;
        RECT  10.490 2.380 11.690 2.780 ;
        RECT  10.495 1.020 11.685 1.420 ;
        RECT  10.250 0.690 10.495 1.420 ;
        RECT  10.250 2.380 10.490 3.380 ;
        RECT  10.245 0.690 10.250 2.780 ;
        RECT  9.350 1.020 10.245 2.780 ;
        RECT  9.050 1.020 9.350 1.420 ;
        RECT  9.050 2.380 9.350 2.780 ;
        RECT  8.810 0.690 9.050 1.420 ;
        RECT  8.810 2.380 9.050 3.380 ;
        RECT  7.610 1.020 8.810 1.420 ;
        RECT  7.610 2.380 8.810 2.780 ;
        RECT  7.370 0.680 7.610 1.420 ;
        RECT  7.370 2.380 7.610 3.380 ;
        END
    END Z
    PIN OE
        ANTENNAGATEAREA 0.7353 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 2.020 5.115 2.755 ;
        RECT  3.885 2.515 4.885 2.755 ;
        RECT  3.645 2.515 3.885 3.225 ;
        RECT  3.150 2.985 3.645 3.225 ;
        RECT  2.920 2.985 3.150 3.455 ;
        RECT  1.760 3.225 2.920 3.455 ;
        RECT  1.530 2.940 1.760 3.455 ;
        RECT  1.030 2.940 1.530 3.170 ;
        RECT  0.980 2.650 1.030 3.170 ;
        RECT  0.800 1.615 0.980 3.170 ;
        RECT  0.650 1.615 0.800 3.030 ;
        END
    END OE
    PIN I
        ANTENNAGATEAREA 1.1574 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 1.595 3.860 1.825 ;
        RECT  2.715 1.595 2.945 2.285 ;
        RECT  1.720 2.055 2.715 2.285 ;
        RECT  1.540 1.585 1.720 2.285 ;
        RECT  1.260 1.585 1.540 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.720 -0.235 12.880 0.235 ;
        RECT  12.340 -0.235 12.720 0.975 ;
        RECT  11.275 -0.235 12.340 0.235 ;
        RECT  10.895 -0.235 11.275 0.790 ;
        RECT  9.835 -0.235 10.895 0.235 ;
        RECT  9.455 -0.235 9.835 0.790 ;
        RECT  8.395 -0.235 9.455 0.235 ;
        RECT  8.015 -0.235 8.395 0.790 ;
        RECT  6.910 -0.235 8.015 0.235 ;
        RECT  6.570 -0.235 6.910 0.715 ;
        RECT  3.420 -0.235 6.570 0.235 ;
        RECT  3.040 -0.235 3.420 0.465 ;
        RECT  1.260 -0.235 3.040 0.235 ;
        RECT  0.880 -0.235 1.260 0.710 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.720 3.685 12.880 4.155 ;
        RECT  12.340 2.570 12.720 4.155 ;
        RECT  11.280 3.685 12.340 4.155 ;
        RECT  10.900 3.030 11.280 4.155 ;
        RECT  9.840 3.685 10.900 4.155 ;
        RECT  9.460 3.030 9.840 4.155 ;
        RECT  8.400 3.685 9.460 4.155 ;
        RECT  8.020 3.030 8.400 4.155 ;
        RECT  6.885 3.685 8.020 4.155 ;
        RECT  6.505 3.015 6.885 4.155 ;
        RECT  5.305 3.685 6.505 4.155 ;
        RECT  4.965 3.455 5.305 4.155 ;
        RECT  3.780 3.685 4.965 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.280 3.685 3.440 4.155 ;
        RECT  0.940 3.440 1.280 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.685 0.690 11.935 1.420 ;
        RECT  11.690 2.380 11.930 3.380 ;
        RECT  10.490 2.380 11.690 2.780 ;
        RECT  10.495 1.020 11.685 1.420 ;
        RECT  10.450 0.690 10.495 1.420 ;
        RECT  10.450 2.380 10.490 3.380 ;
        RECT  9.050 1.020 9.150 1.420 ;
        RECT  9.050 2.380 9.150 2.780 ;
        RECT  8.810 0.690 9.050 1.420 ;
        RECT  8.810 2.380 9.050 3.380 ;
        RECT  7.610 1.020 8.810 1.420 ;
        RECT  7.610 2.380 8.810 2.780 ;
        RECT  7.370 0.680 7.610 1.420 ;
        RECT  7.370 2.380 7.610 3.380 ;
        RECT  7.860 1.880 8.200 2.140 ;
        RECT  6.015 1.910 7.860 2.140 ;
        RECT  6.080 1.430 7.140 1.665 ;
        RECT  5.850 0.465 6.080 1.665 ;
        RECT  5.775 1.910 6.015 3.455 ;
        RECT  4.380 0.465 5.850 0.695 ;
        RECT  5.605 1.910 5.775 2.140 ;
        RECT  4.490 2.985 5.775 3.225 ;
        RECT  5.365 1.020 5.605 2.140 ;
        RECT  5.005 1.020 5.365 1.250 ;
        RECT  4.260 2.985 4.490 3.455 ;
        RECT  4.150 0.465 4.380 2.285 ;
        RECT  4.140 0.935 4.150 2.285 ;
        RECT  2.810 0.935 4.140 1.165 ;
        RECT  3.415 2.055 4.140 2.285 ;
        RECT  3.175 2.055 3.415 2.755 ;
        RECT  2.690 2.515 3.175 2.755 ;
        RECT  2.580 0.465 2.810 1.165 ;
        RECT  2.460 2.515 2.690 2.995 ;
        RECT  1.620 0.465 2.580 0.695 ;
        RECT  2.350 1.485 2.485 1.825 ;
        RECT  2.190 2.765 2.460 2.995 ;
        RECT  2.120 1.105 2.350 1.825 ;
        RECT  0.465 1.105 2.120 1.335 ;
        RECT  0.350 3.225 0.520 3.455 ;
        RECT  0.350 0.465 0.465 1.335 ;
        RECT  0.120 0.465 0.350 3.455 ;
    END
END BUFTD8BWP7T

MACRO CKAN2D0BWP7T
    CLASS CORE ;
    FOREIGN CKAN2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.7440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 0.630 2.660 3.250 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2115 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2034 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.470 0.455 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.830 -0.235 2.800 0.235 ;
        RECT  1.450 -0.235 1.830 0.915 ;
        RECT  0.000 -0.235 1.450 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 3.685 2.800 4.155 ;
        RECT  1.480 3.360 1.735 4.155 ;
        RECT  1.120 3.685 1.480 4.155 ;
        RECT  0.880 3.355 1.120 4.155 ;
        RECT  0.520 3.685 0.880 4.155 ;
        RECT  0.280 3.360 0.520 4.155 ;
        RECT  0.000 3.685 0.280 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.855 1.480 2.085 2.740 ;
        RECT  0.935 2.490 1.855 2.740 ;
        RECT  0.705 0.680 0.935 2.740 ;
        RECT  0.175 0.680 0.705 0.920 ;
    END
END CKAN2D0BWP7T

MACRO CKAN2D1BWP7T
    CLASS CORE ;
    FOREIGN CKAN2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.9096 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 0.610 2.660 3.375 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2520 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2430 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.470 0.455 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.830 -0.235 2.800 0.235 ;
        RECT  1.450 -0.235 1.830 0.880 ;
        RECT  0.000 -0.235 1.450 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 3.685 2.800 4.155 ;
        RECT  1.540 3.095 1.920 4.155 ;
        RECT  0.000 3.685 1.540 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.855 1.480 2.085 2.725 ;
        RECT  0.935 2.475 1.855 2.725 ;
        RECT  0.705 0.650 0.935 2.725 ;
        RECT  0.175 0.650 0.705 0.890 ;
    END
END CKAN2D1BWP7T

MACRO CKAN2D2BWP7T
    CLASS CORE ;
    FOREIGN CKAN2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.0233 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 1.000 3.220 2.710 ;
        RECT  2.970 0.490 2.975 2.710 ;
        RECT  2.940 0.490 2.970 3.410 ;
        RECT  2.725 0.490 2.940 1.240 ;
        RECT  2.730 2.355 2.940 3.410 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.3654 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.570 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3546 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.605 0.455 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 -0.235 3.920 0.235 ;
        RECT  3.380 -0.235 3.760 0.775 ;
        RECT  2.190 -0.235 3.380 0.235 ;
        RECT  1.810 -0.235 2.190 0.720 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.685 3.685 3.920 4.155 ;
        RECT  3.450 2.220 3.685 4.155 ;
        RECT  2.210 3.685 3.450 4.155 ;
        RECT  1.830 2.980 2.210 4.155 ;
        RECT  0.540 3.685 1.830 4.155 ;
        RECT  0.160 2.980 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.255 1.465 2.485 2.725 ;
        RECT  1.290 2.475 2.255 2.725 ;
        RECT  1.060 2.475 1.290 3.375 ;
        RECT  1.010 2.475 1.060 2.725 ;
        RECT  0.780 0.595 1.010 2.725 ;
        RECT  0.245 0.595 0.780 0.835 ;
    END
END CKAN2D2BWP7T

MACRO CKAN2D4BWP7T
    CLASS CORE ;
    FOREIGN CKAN2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.0466 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.440 0.490 5.770 3.205 ;
        RECT  4.870 0.990 5.440 2.550 ;
        RECT  4.255 0.990 4.870 1.340 ;
        RECT  4.255 2.200 4.870 2.550 ;
        RECT  4.005 0.490 4.255 1.340 ;
        RECT  4.000 2.200 4.255 3.205 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.5886 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 1.600 3.040 2.660 ;
        RECT  0.980 2.400 2.760 2.660 ;
        RECT  0.700 1.210 0.980 2.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.5886 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.650 2.230 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 -0.235 6.720 0.235 ;
        RECT  6.110 -0.235 6.490 0.725 ;
        RECT  5.050 -0.235 6.110 0.235 ;
        RECT  4.670 -0.235 5.050 0.720 ;
        RECT  3.555 -0.235 4.670 0.235 ;
        RECT  3.175 -0.235 3.555 0.725 ;
        RECT  0.540 -0.235 3.175 0.235 ;
        RECT  0.160 -0.235 0.540 0.735 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.480 3.685 6.720 4.155 ;
        RECT  6.100 2.305 6.480 4.155 ;
        RECT  5.050 3.685 6.100 4.155 ;
        RECT  4.670 2.780 5.050 4.155 ;
        RECT  3.540 3.685 4.670 4.155 ;
        RECT  3.200 3.450 3.540 4.155 ;
        RECT  2.000 3.685 3.200 4.155 ;
        RECT  1.660 3.450 2.000 4.155 ;
        RECT  0.470 3.685 1.660 4.155 ;
        RECT  0.230 2.360 0.470 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.255 0.990 4.670 1.340 ;
        RECT  4.255 2.200 4.670 2.550 ;
        RECT  4.005 0.490 4.255 1.340 ;
        RECT  4.000 2.200 4.255 3.205 ;
        RECT  3.580 1.610 4.530 1.850 ;
        RECT  3.340 1.140 3.580 3.145 ;
        RECT  2.000 1.140 3.340 1.370 ;
        RECT  0.900 2.900 3.340 3.145 ;
        RECT  0.900 0.465 2.760 0.695 ;
        RECT  1.660 0.965 2.000 1.370 ;
    END
END CKAN2D4BWP7T

MACRO CKAN2D8BWP7T
    CLASS CORE ;
    FOREIGN CKAN2D8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 4.5108 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.610 0.490 9.850 1.305 ;
        RECT  9.610 2.125 9.850 3.260 ;
        RECT  8.410 0.905 9.610 1.305 ;
        RECT  8.410 2.125 9.610 2.525 ;
        RECT  8.170 0.490 8.410 1.305 ;
        RECT  8.170 2.125 8.410 3.260 ;
        RECT  8.010 0.905 8.170 1.305 ;
        RECT  8.010 2.125 8.170 2.525 ;
        RECT  7.110 0.905 8.010 2.525 ;
        RECT  6.970 0.905 7.110 1.280 ;
        RECT  6.970 2.125 7.110 2.525 ;
        RECT  6.730 0.490 6.970 1.280 ;
        RECT  6.730 2.125 6.970 3.260 ;
        RECT  5.560 0.905 6.730 1.280 ;
        RECT  5.530 2.125 6.730 2.525 ;
        RECT  5.280 0.490 5.560 1.280 ;
        RECT  5.290 2.125 5.530 3.260 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 1.1016 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.865 1.670 4.340 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.0746 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.670 2.125 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.200 -0.235 10.080 0.235 ;
        RECT  8.820 -0.235 9.200 0.675 ;
        RECT  7.765 -0.235 8.820 0.235 ;
        RECT  7.385 -0.235 7.765 0.675 ;
        RECT  6.325 -0.235 7.385 0.235 ;
        RECT  5.945 -0.235 6.325 0.675 ;
        RECT  4.875 -0.235 5.945 0.235 ;
        RECT  4.495 -0.235 4.875 0.775 ;
        RECT  3.420 -0.235 4.495 0.235 ;
        RECT  3.040 -0.235 3.420 0.820 ;
        RECT  0.000 -0.235 3.040 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.200 3.685 10.080 4.155 ;
        RECT  8.820 2.775 9.200 4.155 ;
        RECT  7.760 3.685 8.820 4.155 ;
        RECT  7.380 2.775 7.760 4.155 ;
        RECT  6.320 3.685 7.380 4.155 ;
        RECT  5.940 2.775 6.320 4.155 ;
        RECT  4.875 3.685 5.940 4.155 ;
        RECT  4.495 2.960 4.875 4.155 ;
        RECT  3.425 3.685 4.495 4.155 ;
        RECT  3.045 2.960 3.425 4.155 ;
        RECT  1.985 3.685 3.045 4.155 ;
        RECT  1.605 2.960 1.985 4.155 ;
        RECT  0.545 3.685 1.605 4.155 ;
        RECT  0.165 2.960 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.610 0.490 9.850 1.305 ;
        RECT  9.610 2.125 9.850 3.260 ;
        RECT  8.410 0.905 9.610 1.305 ;
        RECT  8.410 2.125 9.610 2.525 ;
        RECT  8.210 0.490 8.410 1.305 ;
        RECT  8.210 2.125 8.410 3.260 ;
        RECT  6.730 0.490 6.910 1.280 ;
        RECT  6.730 2.125 6.910 3.260 ;
        RECT  5.560 0.905 6.730 1.280 ;
        RECT  5.530 2.125 6.730 2.525 ;
        RECT  5.280 0.490 5.560 1.280 ;
        RECT  5.290 2.125 5.530 3.260 ;
        RECT  4.915 1.510 6.840 1.740 ;
        RECT  4.685 1.510 4.915 2.690 ;
        RECT  4.065 2.460 4.685 2.690 ;
        RECT  3.835 0.780 4.065 1.295 ;
        RECT  3.835 2.460 4.065 3.330 ;
        RECT  2.625 1.065 3.835 1.295 ;
        RECT  2.625 2.460 3.835 2.690 ;
        RECT  2.395 0.465 2.625 1.295 ;
        RECT  2.395 2.460 2.625 3.330 ;
        RECT  1.240 0.465 2.395 0.695 ;
        RECT  1.185 2.460 2.395 2.690 ;
        RECT  1.620 0.925 1.960 1.440 ;
        RECT  0.465 1.210 1.620 1.440 ;
        RECT  0.900 0.465 1.240 0.905 ;
        RECT  0.955 2.460 1.185 3.330 ;
        RECT  0.465 2.460 0.955 2.690 ;
        RECT  0.235 0.785 0.465 2.690 ;
    END
END CKAN2D8BWP7T

MACRO CKBD0BWP7T
    CLASS CORE ;
    FOREIGN CKBD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.7440 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 0.485 2.100 3.440 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3042 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.135 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.235 2.240 0.235 ;
        RECT  0.930 -0.235 1.310 0.770 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 3.685 2.240 4.155 ;
        RECT  0.930 2.960 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.260 1.120 1.495 1.795 ;
        RECT  0.470 1.120 1.260 1.350 ;
        RECT  0.345 0.485 0.470 1.350 ;
        RECT  0.345 2.530 0.465 3.420 ;
        RECT  0.115 0.485 0.345 3.420 ;
    END
END CKBD0BWP7T

MACRO CKBD10BWP7T
    CLASS CORE ;
    FOREIGN CKBD10BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 5.6890 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.050 0.470 11.290 1.310 ;
        RECT  11.050 2.135 11.290 3.385 ;
        RECT  9.850 0.910 11.050 1.310 ;
        RECT  9.850 2.135 11.050 2.535 ;
        RECT  9.690 0.540 9.850 1.310 ;
        RECT  9.690 2.135 9.850 3.385 ;
        RECT  9.610 0.540 9.690 3.385 ;
        RECT  8.410 0.910 9.610 2.535 ;
        RECT  8.230 0.540 8.410 3.385 ;
        RECT  8.170 0.540 8.230 1.310 ;
        RECT  8.170 2.135 8.230 3.385 ;
        RECT  6.960 0.910 8.170 1.310 ;
        RECT  6.970 2.135 8.170 2.535 ;
        RECT  6.730 2.135 6.970 3.385 ;
        RECT  6.720 0.475 6.960 1.310 ;
        RECT  5.530 2.135 6.730 2.535 ;
        RECT  5.520 0.910 6.720 1.310 ;
        RECT  5.290 2.135 5.530 3.385 ;
        RECT  5.280 0.475 5.520 1.310 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 1.6920 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 0.760 0.480 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.630 -0.235 11.760 0.235 ;
        RECT  10.250 -0.235 10.630 0.680 ;
        RECT  9.190 -0.235 10.250 0.235 ;
        RECT  8.810 -0.235 9.190 0.680 ;
        RECT  7.760 -0.235 8.810 0.235 ;
        RECT  7.380 -0.235 7.760 0.680 ;
        RECT  6.320 -0.235 7.380 0.235 ;
        RECT  5.940 -0.235 6.320 0.680 ;
        RECT  4.880 -0.235 5.940 0.235 ;
        RECT  4.500 -0.235 4.880 0.830 ;
        RECT  3.430 -0.235 4.500 0.235 ;
        RECT  3.050 -0.235 3.430 0.840 ;
        RECT  1.990 -0.235 3.050 0.235 ;
        RECT  1.610 -0.235 1.990 0.840 ;
        RECT  0.000 -0.235 1.610 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.650 3.685 11.760 4.155 ;
        RECT  10.270 2.765 10.650 4.155 ;
        RECT  9.210 3.685 10.270 4.155 ;
        RECT  8.830 2.765 9.210 4.155 ;
        RECT  7.770 3.685 8.830 4.155 ;
        RECT  7.390 2.765 7.770 4.155 ;
        RECT  6.330 3.685 7.390 4.155 ;
        RECT  5.950 2.765 6.330 4.155 ;
        RECT  4.870 3.685 5.950 4.155 ;
        RECT  4.490 2.580 4.870 4.155 ;
        RECT  3.420 3.685 4.490 4.155 ;
        RECT  3.040 2.580 3.420 4.155 ;
        RECT  1.980 3.685 3.040 4.155 ;
        RECT  1.600 2.580 1.980 4.155 ;
        RECT  0.540 3.685 1.600 4.155 ;
        RECT  0.160 2.580 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.050 0.470 11.290 1.310 ;
        RECT  11.050 2.135 11.290 3.385 ;
        RECT  9.890 0.910 11.050 1.310 ;
        RECT  9.890 2.135 11.050 2.535 ;
        RECT  6.960 0.910 8.030 1.310 ;
        RECT  6.970 2.135 8.030 2.535 ;
        RECT  6.730 2.135 6.970 3.385 ;
        RECT  6.720 0.475 6.960 1.310 ;
        RECT  5.530 2.135 6.730 2.535 ;
        RECT  5.520 0.910 6.720 1.310 ;
        RECT  5.290 2.135 5.530 3.385 ;
        RECT  5.280 0.475 5.520 1.310 ;
        RECT  4.080 1.570 7.695 1.800 ;
        RECT  3.840 0.540 4.080 3.430 ;
        RECT  2.630 1.575 3.840 1.865 ;
        RECT  2.390 0.540 2.630 3.430 ;
        RECT  1.190 1.575 2.390 1.865 ;
        RECT  0.950 0.540 1.190 3.430 ;
    END
END CKBD10BWP7T

MACRO CKBD12BWP7T
    CLASS CORE ;
    FOREIGN CKBD12BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 6.0373 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.770 0.555 12.010 1.310 ;
        RECT  10.570 0.910 11.770 1.310 ;
        RECT  11.050 2.135 11.290 3.365 ;
        RECT  9.850 2.135 11.050 2.535 ;
        RECT  10.330 0.555 10.570 1.310 ;
        RECT  9.690 0.910 10.330 1.310 ;
        RECT  9.690 2.135 9.850 3.380 ;
        RECT  9.610 0.910 9.690 3.380 ;
        RECT  9.130 0.910 9.610 2.535 ;
        RECT  8.890 0.555 9.130 2.535 ;
        RECT  8.410 0.910 8.890 2.535 ;
        RECT  8.230 0.910 8.410 3.380 ;
        RECT  6.960 0.910 8.230 1.310 ;
        RECT  8.170 2.135 8.230 3.380 ;
        RECT  6.970 2.135 8.170 2.535 ;
        RECT  6.730 2.135 6.970 3.380 ;
        RECT  6.720 0.570 6.960 1.310 ;
        RECT  5.530 2.135 6.730 2.535 ;
        RECT  5.520 0.910 6.720 1.310 ;
        RECT  5.290 2.135 5.530 3.380 ;
        RECT  5.280 0.570 5.520 1.310 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 1.9890 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 0.555 0.480 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.350 -0.235 12.320 0.235 ;
        RECT  10.970 -0.235 11.350 0.680 ;
        RECT  9.910 -0.235 10.970 0.235 ;
        RECT  9.530 -0.235 9.910 0.680 ;
        RECT  8.470 -0.235 9.530 0.235 ;
        RECT  8.090 -0.235 8.470 0.680 ;
        RECT  7.760 -0.235 8.090 0.235 ;
        RECT  7.380 -0.235 7.760 0.680 ;
        RECT  6.320 -0.235 7.380 0.235 ;
        RECT  5.940 -0.235 6.320 0.680 ;
        RECT  4.880 -0.235 5.940 0.235 ;
        RECT  4.500 -0.235 4.880 0.755 ;
        RECT  3.430 -0.235 4.500 0.235 ;
        RECT  3.050 -0.235 3.430 0.755 ;
        RECT  1.990 -0.235 3.050 0.235 ;
        RECT  1.610 -0.235 1.990 0.755 ;
        RECT  0.000 -0.235 1.610 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.090 3.685 12.320 4.155 ;
        RECT  11.710 2.520 12.090 4.155 ;
        RECT  10.650 3.685 11.710 4.155 ;
        RECT  10.270 2.765 10.650 4.155 ;
        RECT  9.210 3.685 10.270 4.155 ;
        RECT  8.830 2.765 9.210 4.155 ;
        RECT  7.770 3.685 8.830 4.155 ;
        RECT  7.390 2.765 7.770 4.155 ;
        RECT  6.330 3.685 7.390 4.155 ;
        RECT  5.950 2.765 6.330 4.155 ;
        RECT  4.870 3.685 5.950 4.155 ;
        RECT  4.490 2.495 4.870 4.155 ;
        RECT  3.420 3.685 4.490 4.155 ;
        RECT  3.040 2.490 3.420 4.155 ;
        RECT  1.980 3.685 3.040 4.155 ;
        RECT  1.600 2.495 1.980 4.155 ;
        RECT  0.540 3.685 1.600 4.155 ;
        RECT  0.160 2.545 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.770 0.555 12.010 1.310 ;
        RECT  10.570 0.910 11.770 1.310 ;
        RECT  11.050 2.135 11.290 3.365 ;
        RECT  9.890 2.135 11.050 2.535 ;
        RECT  10.330 0.555 10.570 1.310 ;
        RECT  9.890 0.910 10.330 1.310 ;
        RECT  6.960 0.910 8.030 1.310 ;
        RECT  6.970 2.135 8.030 2.535 ;
        RECT  6.730 2.135 6.970 3.380 ;
        RECT  6.720 0.570 6.960 1.310 ;
        RECT  5.530 2.135 6.730 2.535 ;
        RECT  5.520 0.910 6.720 1.310 ;
        RECT  5.290 2.135 5.530 3.380 ;
        RECT  5.280 0.570 5.520 1.310 ;
        RECT  4.080 1.550 7.690 1.785 ;
        RECT  3.840 0.525 4.080 3.355 ;
        RECT  2.630 1.520 3.840 1.810 ;
        RECT  2.390 0.525 2.630 3.355 ;
        RECT  1.190 1.520 2.390 1.810 ;
        RECT  0.950 0.525 1.190 3.355 ;
    END
END CKBD12BWP7T

MACRO CKBD1BWP7T
    CLASS CORE ;
    FOREIGN CKBD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.9072 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 0.495 2.100 3.405 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3285 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.645 0.980 2.710 ;
        RECT  0.610 1.645 0.700 1.985 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.235 2.240 0.235 ;
        RECT  0.930 -0.235 1.310 0.770 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 3.685 2.240 4.155 ;
        RECT  0.930 3.045 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.290 1.120 1.530 1.460 ;
        RECT  0.470 1.120 1.290 1.350 ;
        RECT  0.370 0.500 0.470 1.350 ;
        RECT  0.370 2.550 0.470 3.450 ;
        RECT  0.140 0.500 0.370 3.450 ;
    END
END CKBD1BWP7T

MACRO CKBD2BWP7T
    CLASS CORE ;
    FOREIGN CKBD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.0233 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.410 1.080 2.660 2.710 ;
        RECT  2.380 0.575 2.410 3.330 ;
        RECT  2.170 0.575 2.380 1.310 ;
        RECT  2.165 2.245 2.380 3.330 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.3717 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 -0.235 3.360 0.235 ;
        RECT  2.820 -0.235 3.200 0.865 ;
        RECT  1.760 -0.235 2.820 0.235 ;
        RECT  1.380 -0.235 1.760 0.815 ;
        RECT  0.000 -0.235 1.380 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 3.685 3.360 4.155 ;
        RECT  2.895 2.250 3.130 4.155 ;
        RECT  1.760 3.685 2.895 4.155 ;
        RECT  1.380 2.295 1.760 4.155 ;
        RECT  0.000 3.685 1.380 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.955 1.540 2.125 1.880 ;
        RECT  0.950 0.525 0.955 1.880 ;
        RECT  0.710 0.525 0.950 3.330 ;
    END
END CKBD2BWP7T

MACRO CKBD3BWP7T
    CLASS CORE ;
    FOREIGN CKBD3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.8730 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.090 2.195 4.195 3.425 ;
        RECT  3.955 1.030 4.090 3.425 ;
        RECT  3.475 1.030 3.955 2.545 ;
        RECT  3.190 0.665 3.475 2.545 ;
        RECT  2.675 2.195 3.190 2.545 ;
        RECT  2.435 2.195 2.675 3.425 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.5544 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.480 1.640 1.230 1.880 ;
        RECT  0.140 0.920 0.480 2.190 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 -0.235 4.480 0.235 ;
        RECT  3.890 -0.235 4.270 0.790 ;
        RECT  2.830 -0.235 3.890 0.235 ;
        RECT  2.450 -0.235 2.830 0.975 ;
        RECT  1.305 -0.235 2.450 0.235 ;
        RECT  0.925 -0.235 1.305 0.945 ;
        RECT  0.000 -0.235 0.925 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 3.685 4.480 4.155 ;
        RECT  3.120 2.775 3.500 4.155 ;
        RECT  2.025 3.685 3.120 4.155 ;
        RECT  1.645 2.650 2.025 4.155 ;
        RECT  0.580 3.685 1.645 4.155 ;
        RECT  0.200 2.630 0.580 4.155 ;
        RECT  0.000 3.685 0.200 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.955 1.710 2.955 1.950 ;
        RECT  1.715 0.635 1.955 2.410 ;
        RECT  1.230 2.150 1.715 2.410 ;
        RECT  0.995 2.150 1.230 3.435 ;
    END
END CKBD3BWP7T

MACRO CKBD4BWP7T
    CLASS CORE ;
    FOREIGN CKBD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.2384 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.555 0.705 4.800 1.545 ;
        RECT  4.090 1.195 4.555 1.545 ;
        RECT  3.840 1.195 4.090 3.430 ;
        RECT  3.360 1.195 3.840 2.590 ;
        RECT  3.190 0.710 3.360 2.590 ;
        RECT  3.115 0.710 3.190 1.545 ;
        RECT  2.630 2.240 3.190 2.590 ;
        RECT  2.390 2.240 2.630 3.430 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.6570 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 0.920 0.480 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.155 -0.235 5.040 0.235 ;
        RECT  3.775 -0.235 4.155 0.955 ;
        RECT  2.710 -0.235 3.775 0.235 ;
        RECT  2.330 -0.235 2.710 0.900 ;
        RECT  1.270 -0.235 2.330 0.235 ;
        RECT  0.890 -0.235 1.270 0.875 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.870 3.685 5.040 4.155 ;
        RECT  4.490 2.300 4.870 4.155 ;
        RECT  3.430 3.685 4.490 4.155 ;
        RECT  3.050 2.915 3.430 4.155 ;
        RECT  1.980 3.685 3.050 4.155 ;
        RECT  1.600 2.300 1.980 4.155 ;
        RECT  0.540 3.685 1.600 4.155 ;
        RECT  0.160 2.470 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.555 0.705 4.800 1.545 ;
        RECT  4.290 1.195 4.555 1.545 ;
        RECT  2.630 2.240 2.990 2.590 ;
        RECT  2.390 2.240 2.630 3.430 ;
        RECT  1.910 1.760 2.910 2.010 ;
        RECT  1.670 0.595 1.910 2.010 ;
        RECT  1.190 1.780 1.670 2.010 ;
        RECT  0.950 1.780 1.190 3.430 ;
    END
END CKBD4BWP7T

MACRO CKBD6BWP7T
    CLASS CORE ;
    FOREIGN CKBD6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 3.2490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.720 0.705 6.965 1.480 ;
        RECT  5.770 1.130 6.720 1.480 ;
        RECT  6.000 2.190 6.250 3.390 ;
        RECT  5.770 2.190 6.000 2.540 ;
        RECT  5.520 1.130 5.770 2.540 ;
        RECT  5.275 0.705 5.520 2.540 ;
        RECT  4.870 1.130 5.275 2.540 ;
        RECT  4.080 1.130 4.870 1.480 ;
        RECT  4.810 2.190 4.870 2.540 ;
        RECT  4.560 2.190 4.810 3.390 ;
        RECT  3.350 2.190 4.560 2.540 ;
        RECT  3.835 0.710 4.080 1.480 ;
        RECT  3.110 2.190 3.350 3.390 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.9990 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.480 1.660 1.445 1.895 ;
        RECT  0.140 0.920 0.480 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.320 -0.235 7.280 0.235 ;
        RECT  5.940 -0.235 6.320 0.900 ;
        RECT  4.875 -0.235 5.940 0.235 ;
        RECT  4.495 -0.235 4.875 0.900 ;
        RECT  3.430 -0.235 4.495 0.235 ;
        RECT  3.050 -0.235 3.430 1.005 ;
        RECT  2.710 -0.235 3.050 0.235 ;
        RECT  2.330 -0.235 2.710 1.020 ;
        RECT  1.270 -0.235 2.330 0.235 ;
        RECT  0.890 -0.235 1.270 0.995 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.035 3.685 7.280 4.155 ;
        RECT  6.655 2.300 7.035 4.155 ;
        RECT  5.590 3.685 6.655 4.155 ;
        RECT  5.210 2.770 5.590 4.155 ;
        RECT  4.145 3.685 5.210 4.155 ;
        RECT  3.765 2.770 4.145 4.155 ;
        RECT  2.700 3.685 3.765 4.155 ;
        RECT  2.320 2.300 2.700 4.155 ;
        RECT  1.260 3.685 2.320 4.155 ;
        RECT  0.880 2.975 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.720 0.705 6.965 1.480 ;
        RECT  5.970 1.130 6.720 1.480 ;
        RECT  6.000 2.190 6.250 3.390 ;
        RECT  5.970 2.190 6.000 2.540 ;
        RECT  4.080 1.130 4.670 1.480 ;
        RECT  4.560 2.190 4.670 3.390 ;
        RECT  3.350 2.190 4.560 2.540 ;
        RECT  3.835 0.710 4.080 1.480 ;
        RECT  3.110 2.190 3.350 3.390 ;
        RECT  1.910 1.710 4.570 1.960 ;
        RECT  1.675 0.740 1.910 3.390 ;
        RECT  1.670 2.440 1.675 3.390 ;
        RECT  0.470 2.440 1.670 2.685 ;
        RECT  0.230 2.440 0.470 3.385 ;
    END
END CKBD6BWP7T

MACRO CKBD8BWP7T
    CLASS CORE ;
    FOREIGN CKBD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 3.9044 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.165 2.245 8.415 3.340 ;
        RECT  6.970 2.245 8.165 2.645 ;
        RECT  7.440 0.655 7.685 1.500 ;
        RECT  6.890 1.100 7.440 1.500 ;
        RECT  6.890 2.245 6.970 3.340 ;
        RECT  6.720 1.100 6.890 3.340 ;
        RECT  6.240 1.100 6.720 2.645 ;
        RECT  5.995 0.655 6.240 2.645 ;
        RECT  5.990 1.100 5.995 2.645 ;
        RECT  4.800 1.100 5.990 1.500 ;
        RECT  5.530 2.245 5.990 2.645 ;
        RECT  5.280 2.245 5.530 3.340 ;
        RECT  4.070 2.245 5.280 2.645 ;
        RECT  4.555 0.660 4.800 1.500 ;
        RECT  3.830 2.245 4.070 3.340 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 1.2186 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.480 1.660 1.915 1.895 ;
        RECT  0.140 0.920 0.480 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.480 -0.235 8.960 0.235 ;
        RECT  8.100 -0.235 8.480 1.005 ;
        RECT  7.040 -0.235 8.100 0.235 ;
        RECT  6.660 -0.235 7.040 0.870 ;
        RECT  5.595 -0.235 6.660 0.235 ;
        RECT  5.215 -0.235 5.595 0.870 ;
        RECT  4.150 -0.235 5.215 0.235 ;
        RECT  3.770 -0.235 4.150 1.005 ;
        RECT  3.430 -0.235 3.770 0.235 ;
        RECT  3.050 -0.235 3.430 0.970 ;
        RECT  1.990 -0.235 3.050 0.235 ;
        RECT  1.610 -0.235 1.990 0.920 ;
        RECT  0.000 -0.235 1.610 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.755 3.685 8.960 4.155 ;
        RECT  7.375 2.920 7.755 4.155 ;
        RECT  6.310 3.685 7.375 4.155 ;
        RECT  5.930 2.920 6.310 4.155 ;
        RECT  4.865 3.685 5.930 4.155 ;
        RECT  4.485 2.920 4.865 4.155 ;
        RECT  3.420 3.685 4.485 4.155 ;
        RECT  3.040 2.300 3.420 4.155 ;
        RECT  1.980 3.685 3.040 4.155 ;
        RECT  1.600 2.745 1.980 4.155 ;
        RECT  0.540 3.685 1.600 4.155 ;
        RECT  0.160 2.725 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.165 2.245 8.415 3.340 ;
        RECT  7.090 2.245 8.165 2.645 ;
        RECT  7.440 0.655 7.685 1.500 ;
        RECT  7.090 1.100 7.440 1.500 ;
        RECT  4.800 1.100 5.790 1.500 ;
        RECT  5.530 2.245 5.790 2.645 ;
        RECT  5.280 2.245 5.530 3.340 ;
        RECT  4.070 2.245 5.280 2.645 ;
        RECT  4.555 0.660 4.800 1.500 ;
        RECT  3.830 2.245 4.070 3.340 ;
        RECT  2.630 1.730 5.290 1.980 ;
        RECT  2.395 0.620 2.630 3.340 ;
        RECT  1.190 1.150 2.395 1.385 ;
        RECT  1.190 2.245 2.395 2.480 ;
        RECT  0.955 0.620 1.190 1.385 ;
        RECT  0.955 2.245 1.190 3.435 ;
    END
END CKBD8BWP7T

MACRO CKLHQD1BWP7T
    CLASS CORE ;
    FOREIGN CKLHQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.0896 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.715 0.495 11.060 3.235 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 1.680 1.540 2.710 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.5355 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.660 7.140 2.710 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.240 -0.235 11.200 0.235 ;
        RECT  9.995 -0.235 10.240 1.250 ;
        RECT  9.585 -0.235 9.995 0.235 ;
        RECT  9.245 -0.235 9.585 0.470 ;
        RECT  5.515 -0.235 9.245 0.235 ;
        RECT  5.175 -0.235 5.515 0.465 ;
        RECT  3.915 -0.235 5.175 0.235 ;
        RECT  3.685 -0.235 3.915 0.840 ;
        RECT  1.105 -0.235 3.685 0.235 ;
        RECT  0.725 -0.235 1.105 1.265 ;
        RECT  0.000 -0.235 0.725 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.175 3.685 11.200 4.155 ;
        RECT  9.835 3.450 10.175 4.155 ;
        RECT  8.875 3.685 9.835 4.155 ;
        RECT  8.535 3.450 8.875 4.155 ;
        RECT  5.990 3.685 8.535 4.155 ;
        RECT  5.610 3.055 5.990 4.155 ;
        RECT  3.615 3.685 5.610 4.155 ;
        RECT  3.385 3.135 3.615 4.155 ;
        RECT  0.540 3.685 3.385 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.195 1.600 10.430 3.220 ;
        RECT  7.675 2.980 10.195 3.220 ;
        RECT  9.525 0.975 9.765 2.655 ;
        RECT  9.215 0.975 9.525 1.205 ;
        RECT  8.330 2.425 9.525 2.655 ;
        RECT  8.855 1.710 9.225 1.945 ;
        RECT  8.615 0.465 8.855 1.945 ;
        RECT  6.055 0.465 8.615 0.705 ;
        RECT  8.085 1.640 8.330 2.655 ;
        RECT  7.675 1.015 8.120 1.255 ;
        RECT  7.435 1.015 7.675 3.220 ;
        RECT  7.055 2.980 7.435 3.220 ;
        RECT  6.595 1.010 6.715 1.255 ;
        RECT  6.595 3.190 6.695 3.420 ;
        RECT  6.355 1.010 6.595 3.420 ;
        RECT  6.315 1.980 6.355 3.420 ;
        RECT  5.450 1.980 6.315 2.320 ;
        RECT  5.815 0.465 6.055 0.925 ;
        RECT  4.640 0.695 5.815 0.925 ;
        RECT  5.200 1.170 5.375 1.420 ;
        RECT  4.970 1.170 5.200 3.455 ;
        RECT  4.075 3.225 4.970 3.455 ;
        RECT  4.630 0.500 4.640 0.925 ;
        RECT  4.545 0.500 4.630 2.230 ;
        RECT  4.390 0.500 4.545 2.805 ;
        RECT  4.305 2.000 4.390 2.805 ;
        RECT  3.100 2.000 4.305 2.230 ;
        RECT  2.695 1.500 4.160 1.740 ;
        RECT  3.845 2.675 4.075 3.455 ;
        RECT  3.115 2.675 3.845 2.905 ;
        RECT  2.885 2.675 3.115 3.275 ;
        RECT  2.045 0.465 2.990 0.695 ;
        RECT  2.360 3.035 2.885 3.275 ;
        RECT  2.655 0.930 2.695 1.740 ;
        RECT  2.425 0.930 2.655 2.750 ;
        RECT  2.015 2.520 2.425 2.750 ;
        RECT  1.815 0.465 2.045 2.220 ;
    END
END CKLHQD1BWP7T

MACRO CKLHQD2BWP7T
    CLASS CORE ;
    FOREIGN CKLHQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.1445 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.810 1.210 11.060 2.710 ;
        RECT  10.805 0.490 10.810 2.710 ;
        RECT  10.780 0.490 10.805 3.345 ;
        RECT  10.565 0.490 10.780 1.465 ;
        RECT  10.565 2.465 10.780 3.345 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 1.680 1.540 2.710 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.5355 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.660 7.140 2.710 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.535 -0.235 11.760 0.235 ;
        RECT  11.290 -0.235 11.535 1.305 ;
        RECT  10.090 -0.235 11.290 0.235 ;
        RECT  9.845 -0.235 10.090 1.305 ;
        RECT  9.465 -0.235 9.845 0.235 ;
        RECT  9.095 -0.235 9.465 0.470 ;
        RECT  5.515 -0.235 9.095 0.235 ;
        RECT  5.175 -0.235 5.515 0.465 ;
        RECT  3.915 -0.235 5.175 0.235 ;
        RECT  3.685 -0.235 3.915 0.840 ;
        RECT  1.105 -0.235 3.685 0.235 ;
        RECT  0.725 -0.235 1.105 1.265 ;
        RECT  0.000 -0.235 0.725 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.530 3.685 11.760 4.155 ;
        RECT  11.295 2.685 11.530 4.155 ;
        RECT  10.095 3.685 11.295 4.155 ;
        RECT  9.755 3.245 10.095 4.155 ;
        RECT  8.595 3.685 9.755 4.155 ;
        RECT  8.255 3.450 8.595 4.155 ;
        RECT  5.990 3.685 8.255 4.155 ;
        RECT  5.610 3.055 5.990 4.155 ;
        RECT  3.615 3.685 5.610 4.155 ;
        RECT  3.385 3.135 3.615 4.155 ;
        RECT  0.540 3.685 3.385 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.045 1.600 10.280 3.000 ;
        RECT  7.675 2.760 10.045 3.000 ;
        RECT  9.385 0.975 9.615 2.530 ;
        RECT  9.055 0.975 9.385 1.205 ;
        RECT  8.270 2.300 9.385 2.530 ;
        RECT  8.780 1.710 9.155 1.945 ;
        RECT  8.540 0.465 8.780 1.945 ;
        RECT  6.055 0.465 8.540 0.705 ;
        RECT  8.025 1.640 8.270 2.530 ;
        RECT  7.675 1.015 8.060 1.255 ;
        RECT  7.435 1.015 7.675 3.220 ;
        RECT  7.055 2.980 7.435 3.220 ;
        RECT  6.595 1.010 6.715 1.255 ;
        RECT  6.595 3.190 6.695 3.420 ;
        RECT  6.355 1.010 6.595 3.420 ;
        RECT  6.315 1.980 6.355 3.420 ;
        RECT  5.450 1.980 6.315 2.320 ;
        RECT  5.815 0.465 6.055 0.925 ;
        RECT  4.640 0.695 5.815 0.925 ;
        RECT  5.200 1.170 5.375 1.420 ;
        RECT  4.970 1.170 5.200 3.455 ;
        RECT  4.075 3.225 4.970 3.455 ;
        RECT  4.630 0.500 4.640 0.925 ;
        RECT  4.545 0.500 4.630 2.230 ;
        RECT  4.390 0.500 4.545 2.805 ;
        RECT  4.305 2.000 4.390 2.805 ;
        RECT  3.100 2.000 4.305 2.230 ;
        RECT  2.695 1.500 4.160 1.740 ;
        RECT  3.845 2.675 4.075 3.455 ;
        RECT  3.115 2.675 3.845 2.905 ;
        RECT  2.885 2.675 3.115 3.275 ;
        RECT  2.045 0.465 2.990 0.695 ;
        RECT  2.360 3.035 2.885 3.275 ;
        RECT  2.655 0.930 2.695 1.740 ;
        RECT  2.425 0.930 2.655 2.750 ;
        RECT  2.015 2.520 2.425 2.750 ;
        RECT  1.815 0.465 2.045 2.220 ;
    END
END CKLHQD2BWP7T

MACRO CKLHQD4BWP7T
    CLASS CORE ;
    FOREIGN CKLHQD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 2.1384 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.815 0.495 13.050 3.455 ;
        RECT  12.810 1.020 12.815 3.455 ;
        RECT  12.150 1.020 12.810 2.530 ;
        RECT  11.610 1.020 12.150 1.370 ;
        RECT  11.610 2.180 12.150 2.530 ;
        RECT  11.370 0.485 11.610 1.370 ;
        RECT  11.370 2.180 11.610 3.455 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 1.680 1.540 2.710 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.8685 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.160 1.820 9.755 2.050 ;
        RECT  8.930 1.820 9.160 2.525 ;
        RECT  7.445 2.295 8.930 2.525 ;
        RECT  7.215 1.820 7.445 2.525 ;
        RECT  6.180 1.820 7.215 2.100 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.765 -0.235 14.000 0.235 ;
        RECT  13.535 -0.235 13.765 1.275 ;
        RECT  12.400 -0.235 13.535 0.235 ;
        RECT  12.020 -0.235 12.400 0.790 ;
        RECT  10.960 -0.235 12.020 0.235 ;
        RECT  10.580 -0.235 10.960 0.670 ;
        RECT  9.520 -0.235 10.580 0.235 ;
        RECT  9.140 -0.235 9.520 0.670 ;
        RECT  8.060 -0.235 9.140 0.235 ;
        RECT  7.720 -0.235 8.060 0.740 ;
        RECT  5.505 -0.235 7.720 0.235 ;
        RECT  5.165 -0.235 5.505 0.465 ;
        RECT  3.915 -0.235 5.165 0.235 ;
        RECT  3.685 -0.235 3.915 0.725 ;
        RECT  1.105 -0.235 3.685 0.235 ;
        RECT  0.725 -0.235 1.105 1.265 ;
        RECT  0.000 -0.235 0.725 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.765 3.685 14.000 4.155 ;
        RECT  13.535 2.670 13.765 4.155 ;
        RECT  12.400 3.685 13.535 4.155 ;
        RECT  12.020 2.775 12.400 4.155 ;
        RECT  10.860 3.685 12.020 4.155 ;
        RECT  10.520 3.455 10.860 4.155 ;
        RECT  8.180 3.685 10.520 4.155 ;
        RECT  7.800 3.245 8.180 4.155 ;
        RECT  5.985 3.685 7.800 4.155 ;
        RECT  5.605 3.055 5.985 4.155 ;
        RECT  3.615 3.685 5.605 4.155 ;
        RECT  3.385 3.135 3.615 4.155 ;
        RECT  0.540 3.685 3.385 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.610 1.020 11.950 1.370 ;
        RECT  11.610 2.180 11.950 2.530 ;
        RECT  11.370 0.485 11.610 1.370 ;
        RECT  11.370 2.180 11.610 3.455 ;
        RECT  10.890 1.655 11.840 1.900 ;
        RECT  10.650 0.900 10.890 3.225 ;
        RECT  10.220 0.900 10.650 1.130 ;
        RECT  10.250 2.985 10.650 3.225 ;
        RECT  10.165 1.360 10.395 2.610 ;
        RECT  10.010 2.985 10.250 3.455 ;
        RECT  9.880 0.465 10.220 1.130 ;
        RECT  8.400 1.360 10.165 1.590 ;
        RECT  9.780 2.380 10.165 2.610 ;
        RECT  9.160 3.215 10.010 3.455 ;
        RECT  8.780 0.900 9.880 1.130 ;
        RECT  9.550 2.380 9.780 2.985 ;
        RECT  7.035 2.755 9.550 2.985 ;
        RECT  8.440 0.465 8.780 1.130 ;
        RECT  8.170 1.360 8.400 2.000 ;
        RECT  7.990 1.360 8.170 1.615 ;
        RECT  7.760 1.015 7.990 1.615 ;
        RECT  7.000 1.015 7.760 1.255 ;
        RECT  5.975 0.465 6.980 0.695 ;
        RECT  6.405 2.505 6.635 3.360 ;
        RECT  6.345 0.965 6.575 1.385 ;
        RECT  5.665 2.505 6.405 2.735 ;
        RECT  5.895 1.155 6.345 1.385 ;
        RECT  5.735 0.465 5.975 0.925 ;
        RECT  5.665 1.155 5.895 1.865 ;
        RECT  4.690 0.695 5.735 0.925 ;
        RECT  5.435 1.635 5.665 2.735 ;
        RECT  5.110 1.170 5.310 1.420 ;
        RECT  5.110 3.080 5.195 3.455 ;
        RECT  4.880 1.170 5.110 3.455 ;
        RECT  4.075 3.225 4.880 3.455 ;
        RECT  4.630 0.465 4.690 0.925 ;
        RECT  4.540 0.465 4.630 2.230 ;
        RECT  4.390 0.465 4.540 2.805 ;
        RECT  4.350 0.465 4.390 0.695 ;
        RECT  4.305 2.000 4.390 2.805 ;
        RECT  3.100 2.000 4.305 2.230 ;
        RECT  2.695 1.500 4.160 1.740 ;
        RECT  3.845 2.675 4.075 3.455 ;
        RECT  3.115 2.675 3.845 2.905 ;
        RECT  2.885 2.675 3.115 3.275 ;
        RECT  2.045 0.465 2.990 0.695 ;
        RECT  2.360 3.035 2.885 3.275 ;
        RECT  2.655 0.930 2.695 1.740 ;
        RECT  2.425 0.930 2.655 2.750 ;
        RECT  2.015 2.520 2.425 2.750 ;
        RECT  1.815 0.465 2.045 2.220 ;
    END
END CKLHQD4BWP7T

MACRO CKLHQD6BWP7T
    CLASS CORE ;
    FOREIGN CKLHQD6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 3.0780 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.495 0.495 14.730 1.370 ;
        RECT  14.490 2.180 14.730 3.110 ;
        RECT  14.170 1.020 14.495 1.370 ;
        RECT  14.170 2.180 14.490 2.530 ;
        RECT  13.290 1.020 14.170 2.530 ;
        RECT  13.270 0.495 13.290 3.110 ;
        RECT  13.055 0.495 13.270 1.370 ;
        RECT  13.050 2.180 13.270 3.110 ;
        RECT  11.850 1.020 13.055 1.370 ;
        RECT  11.850 2.180 13.050 2.530 ;
        RECT  11.610 0.495 11.850 1.370 ;
        RECT  11.610 2.180 11.850 3.110 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 1.680 1.540 2.710 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.8829 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.160 1.780 9.755 2.010 ;
        RECT  8.930 1.780 9.160 2.525 ;
        RECT  7.700 2.295 8.930 2.525 ;
        RECT  7.105 1.770 7.700 2.525 ;
        RECT  6.860 1.600 7.105 2.525 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.520 -0.235 15.680 0.235 ;
        RECT  15.140 -0.235 15.520 1.255 ;
        RECT  14.080 -0.235 15.140 0.235 ;
        RECT  13.700 -0.235 14.080 0.790 ;
        RECT  12.640 -0.235 13.700 0.235 ;
        RECT  12.260 -0.235 12.640 0.790 ;
        RECT  11.160 -0.235 12.260 0.235 ;
        RECT  10.780 -0.235 11.160 0.560 ;
        RECT  9.640 -0.235 10.780 0.235 ;
        RECT  9.260 -0.235 9.640 0.560 ;
        RECT  8.100 -0.235 9.260 0.235 ;
        RECT  7.760 -0.235 8.100 0.555 ;
        RECT  5.505 -0.235 7.760 0.235 ;
        RECT  5.165 -0.235 5.505 0.465 ;
        RECT  3.915 -0.235 5.165 0.235 ;
        RECT  3.685 -0.235 3.915 0.725 ;
        RECT  1.105 -0.235 3.685 0.235 ;
        RECT  0.725 -0.235 1.105 1.265 ;
        RECT  0.000 -0.235 0.725 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.520 3.685 15.680 4.155 ;
        RECT  15.140 2.300 15.520 4.155 ;
        RECT  14.080 3.685 15.140 4.155 ;
        RECT  13.700 2.775 14.080 4.155 ;
        RECT  12.640 3.685 13.700 4.155 ;
        RECT  12.260 2.775 12.640 4.155 ;
        RECT  11.005 3.685 12.260 4.155 ;
        RECT  10.665 3.455 11.005 4.155 ;
        RECT  8.180 3.685 10.665 4.155 ;
        RECT  7.800 3.245 8.180 4.155 ;
        RECT  5.985 3.685 7.800 4.155 ;
        RECT  5.605 3.055 5.985 4.155 ;
        RECT  3.615 3.685 5.605 4.155 ;
        RECT  3.385 3.135 3.615 4.155 ;
        RECT  0.540 3.685 3.385 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.495 0.495 14.730 1.370 ;
        RECT  14.490 2.180 14.730 3.110 ;
        RECT  14.370 1.020 14.495 1.370 ;
        RECT  14.370 2.180 14.490 2.530 ;
        RECT  13.055 0.495 13.070 1.370 ;
        RECT  13.050 2.180 13.070 3.110 ;
        RECT  11.850 1.020 13.055 1.370 ;
        RECT  11.850 2.180 13.050 2.530 ;
        RECT  11.610 0.495 11.850 1.370 ;
        RECT  11.610 2.180 11.850 3.110 ;
        RECT  11.130 1.655 13.020 1.900 ;
        RECT  10.890 0.860 11.130 3.225 ;
        RECT  10.380 0.860 10.890 1.090 ;
        RECT  10.250 2.985 10.890 3.225 ;
        RECT  10.325 1.320 10.555 2.610 ;
        RECT  10.040 0.465 10.380 1.090 ;
        RECT  8.400 1.320 10.325 1.550 ;
        RECT  9.780 2.380 10.325 2.610 ;
        RECT  10.010 2.985 10.250 3.455 ;
        RECT  8.860 0.860 10.040 1.090 ;
        RECT  9.160 3.215 10.010 3.455 ;
        RECT  9.550 2.380 9.780 2.985 ;
        RECT  7.335 2.755 9.550 2.985 ;
        RECT  8.520 0.465 8.860 1.090 ;
        RECT  8.180 1.320 8.400 2.000 ;
        RECT  8.170 1.015 8.180 2.000 ;
        RECT  7.950 1.015 8.170 1.615 ;
        RECT  7.000 1.015 7.950 1.255 ;
        RECT  7.105 2.755 7.335 3.375 ;
        RECT  5.975 0.465 6.980 0.695 ;
        RECT  6.575 3.190 6.690 3.420 ;
        RECT  6.345 0.965 6.575 3.420 ;
        RECT  5.435 1.980 6.345 2.320 ;
        RECT  5.735 0.465 5.975 0.925 ;
        RECT  4.690 0.695 5.735 0.925 ;
        RECT  5.110 1.170 5.310 1.420 ;
        RECT  5.110 3.080 5.195 3.455 ;
        RECT  4.880 1.170 5.110 3.455 ;
        RECT  4.075 3.225 4.880 3.455 ;
        RECT  4.630 0.465 4.690 0.925 ;
        RECT  4.540 0.465 4.630 2.230 ;
        RECT  4.390 0.465 4.540 2.805 ;
        RECT  4.350 0.465 4.390 0.695 ;
        RECT  4.305 2.000 4.390 2.805 ;
        RECT  3.100 2.000 4.305 2.230 ;
        RECT  2.695 1.500 4.160 1.740 ;
        RECT  3.845 2.675 4.075 3.455 ;
        RECT  3.115 2.675 3.845 2.905 ;
        RECT  2.885 2.675 3.115 3.275 ;
        RECT  2.045 0.465 2.990 0.695 ;
        RECT  2.360 3.035 2.885 3.275 ;
        RECT  2.655 0.930 2.695 1.740 ;
        RECT  2.425 0.930 2.655 2.750 ;
        RECT  2.015 2.520 2.425 2.750 ;
        RECT  1.815 0.465 2.045 2.220 ;
    END
END CKLHQD6BWP7T

MACRO CKLHQD8BWP7T
    CLASS CORE ;
    FOREIGN CKLHQD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 4.3008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.175 0.485 16.410 1.370 ;
        RECT  16.170 2.180 16.410 3.135 ;
        RECT  15.290 1.020 16.175 1.370 ;
        RECT  15.290 2.180 16.170 2.530 ;
        RECT  14.970 1.020 15.290 2.530 ;
        RECT  14.735 0.485 14.970 3.135 ;
        RECT  14.730 1.020 14.735 3.135 ;
        RECT  14.390 1.020 14.730 2.530 ;
        RECT  13.530 1.020 14.390 1.370 ;
        RECT  13.530 2.180 14.390 2.530 ;
        RECT  13.295 0.485 13.530 1.370 ;
        RECT  13.290 2.180 13.530 3.135 ;
        RECT  12.090 1.020 13.295 1.370 ;
        RECT  12.090 2.180 13.290 2.530 ;
        RECT  11.850 0.485 12.090 1.370 ;
        RECT  11.850 2.180 12.090 3.135 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3222 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.145 1.680 1.540 2.710 ;
        END
    END E
    PIN CPN
        ANTENNAGATEAREA 0.8829 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.320 1.780 9.915 2.010 ;
        RECT  9.090 1.780 9.320 2.525 ;
        RECT  7.700 2.295 9.090 2.525 ;
        RECT  7.105 1.770 7.700 2.525 ;
        RECT  6.860 1.600 7.105 2.525 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.200 -0.235 17.360 0.235 ;
        RECT  16.820 -0.235 17.200 1.225 ;
        RECT  15.760 -0.235 16.820 0.235 ;
        RECT  15.380 -0.235 15.760 0.790 ;
        RECT  14.320 -0.235 15.380 0.235 ;
        RECT  13.940 -0.235 14.320 0.790 ;
        RECT  12.880 -0.235 13.940 0.235 ;
        RECT  12.500 -0.235 12.880 0.790 ;
        RECT  11.320 -0.235 12.500 0.235 ;
        RECT  10.940 -0.235 11.320 0.560 ;
        RECT  9.800 -0.235 10.940 0.235 ;
        RECT  9.420 -0.235 9.800 0.560 ;
        RECT  8.260 -0.235 9.420 0.235 ;
        RECT  7.920 -0.235 8.260 0.555 ;
        RECT  5.505 -0.235 7.920 0.235 ;
        RECT  5.165 -0.235 5.505 0.465 ;
        RECT  3.915 -0.235 5.165 0.235 ;
        RECT  3.685 -0.235 3.915 0.725 ;
        RECT  1.105 -0.235 3.685 0.235 ;
        RECT  0.725 -0.235 1.105 1.265 ;
        RECT  0.000 -0.235 0.725 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.200 3.685 17.360 4.155 ;
        RECT  16.820 2.300 17.200 4.155 ;
        RECT  15.760 3.685 16.820 4.155 ;
        RECT  15.380 2.775 15.760 4.155 ;
        RECT  14.320 3.685 15.380 4.155 ;
        RECT  13.940 2.775 14.320 4.155 ;
        RECT  12.880 3.685 13.940 4.155 ;
        RECT  12.500 2.775 12.880 4.155 ;
        RECT  11.165 3.685 12.500 4.155 ;
        RECT  10.825 3.455 11.165 4.155 ;
        RECT  8.340 3.685 10.825 4.155 ;
        RECT  7.960 3.245 8.340 4.155 ;
        RECT  5.985 3.685 7.960 4.155 ;
        RECT  5.605 3.055 5.985 4.155 ;
        RECT  3.615 3.685 5.605 4.155 ;
        RECT  3.385 3.135 3.615 4.155 ;
        RECT  0.540 3.685 3.385 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.175 0.485 16.410 1.370 ;
        RECT  16.170 2.180 16.410 3.135 ;
        RECT  15.490 1.020 16.175 1.370 ;
        RECT  15.490 2.180 16.170 2.530 ;
        RECT  13.530 1.020 14.190 1.370 ;
        RECT  13.530 2.180 14.190 2.530 ;
        RECT  13.295 0.485 13.530 1.370 ;
        RECT  13.290 2.180 13.530 3.135 ;
        RECT  12.090 1.020 13.295 1.370 ;
        RECT  12.090 2.180 13.290 2.530 ;
        RECT  11.850 0.485 12.090 1.370 ;
        RECT  11.850 2.180 12.090 3.135 ;
        RECT  11.290 1.655 13.650 1.900 ;
        RECT  11.050 0.860 11.290 3.225 ;
        RECT  10.540 0.860 11.050 1.090 ;
        RECT  10.410 2.985 11.050 3.225 ;
        RECT  10.485 1.320 10.715 2.610 ;
        RECT  10.200 0.465 10.540 1.090 ;
        RECT  8.560 1.320 10.485 1.550 ;
        RECT  9.940 2.380 10.485 2.610 ;
        RECT  10.170 2.985 10.410 3.455 ;
        RECT  9.020 0.860 10.200 1.090 ;
        RECT  9.320 3.215 10.170 3.455 ;
        RECT  9.710 2.380 9.940 2.985 ;
        RECT  7.335 2.755 9.710 2.985 ;
        RECT  8.680 0.465 9.020 1.090 ;
        RECT  8.340 1.320 8.560 2.000 ;
        RECT  8.330 1.015 8.340 2.000 ;
        RECT  8.110 1.015 8.330 1.615 ;
        RECT  7.160 1.015 8.110 1.255 ;
        RECT  7.105 2.755 7.335 3.375 ;
        RECT  5.975 0.465 6.980 0.695 ;
        RECT  6.575 3.190 6.690 3.420 ;
        RECT  6.345 0.965 6.575 3.420 ;
        RECT  5.435 1.980 6.345 2.320 ;
        RECT  5.735 0.465 5.975 0.925 ;
        RECT  4.690 0.695 5.735 0.925 ;
        RECT  5.110 1.170 5.310 1.420 ;
        RECT  5.110 3.080 5.195 3.455 ;
        RECT  4.880 1.170 5.110 3.455 ;
        RECT  4.075 3.225 4.880 3.455 ;
        RECT  4.630 0.465 4.690 0.925 ;
        RECT  4.540 0.465 4.630 2.230 ;
        RECT  4.390 0.465 4.540 2.805 ;
        RECT  4.350 0.465 4.390 0.695 ;
        RECT  4.305 2.000 4.390 2.805 ;
        RECT  3.100 2.000 4.305 2.230 ;
        RECT  2.695 1.500 4.160 1.740 ;
        RECT  3.845 2.675 4.075 3.455 ;
        RECT  3.115 2.675 3.845 2.905 ;
        RECT  2.885 2.675 3.115 3.275 ;
        RECT  2.045 0.465 2.990 0.695 ;
        RECT  2.360 3.035 2.885 3.275 ;
        RECT  2.655 0.930 2.695 1.740 ;
        RECT  2.425 0.930 2.655 2.750 ;
        RECT  2.015 2.520 2.425 2.750 ;
        RECT  1.815 0.465 2.045 2.220 ;
    END
END CKLHQD8BWP7T

MACRO CKLNQD1BWP7T
    CLASS CORE ;
    FOREIGN CKLNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 0.9096 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.050 0.860 9.380 3.195 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.680 1.555 2.710 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.4653 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.660 7.140 2.710 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.570 -0.235 9.520 0.235 ;
        RECT  8.330 -0.235 8.570 1.190 ;
        RECT  5.515 -0.235 8.330 0.235 ;
        RECT  5.175 -0.235 5.515 0.465 ;
        RECT  3.885 -0.235 5.175 0.235 ;
        RECT  3.655 -0.235 3.885 0.860 ;
        RECT  1.265 -0.235 3.655 0.235 ;
        RECT  0.885 -0.235 1.265 0.820 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.635 3.685 9.520 4.155 ;
        RECT  8.255 3.030 8.635 4.155 ;
        RECT  7.140 3.685 8.255 4.155 ;
        RECT  6.800 3.450 7.140 4.155 ;
        RECT  5.895 3.685 6.800 4.155 ;
        RECT  5.515 2.870 5.895 4.155 ;
        RECT  3.615 3.685 5.515 4.155 ;
        RECT  3.380 2.995 3.615 4.155 ;
        RECT  0.540 3.685 3.380 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.535 1.600 8.765 2.800 ;
        RECT  7.850 2.560 8.535 2.800 ;
        RECT  7.850 0.465 8.090 2.330 ;
        RECT  6.055 0.465 7.850 0.705 ;
        RECT  7.610 2.560 7.850 3.335 ;
        RECT  7.600 2.560 7.610 2.800 ;
        RECT  7.370 0.935 7.600 2.800 ;
        RECT  7.130 0.935 7.370 1.175 ;
        RECT  6.595 0.935 6.715 1.180 ;
        RECT  6.365 0.935 6.595 3.050 ;
        RECT  6.315 2.030 6.365 3.050 ;
        RECT  5.315 2.030 6.315 2.270 ;
        RECT  5.815 0.465 6.055 0.925 ;
        RECT  4.610 0.695 5.815 0.925 ;
        RECT  5.085 1.170 5.375 1.420 ;
        RECT  4.830 1.170 5.085 3.455 ;
        RECT  4.075 3.225 4.830 3.455 ;
        RECT  4.600 0.515 4.610 0.925 ;
        RECT  4.370 0.515 4.600 2.760 ;
        RECT  4.310 1.995 4.370 2.760 ;
        RECT  3.425 1.995 4.310 2.225 ;
        RECT  3.425 1.235 4.125 1.575 ;
        RECT  3.845 2.495 4.075 3.455 ;
        RECT  2.965 2.495 3.845 2.725 ;
        RECT  3.195 0.570 3.425 1.575 ;
        RECT  3.195 1.855 3.425 2.225 ;
        RECT  2.430 0.570 3.195 0.805 ;
        RECT  2.735 1.115 2.965 3.455 ;
        RECT  1.850 3.215 2.735 3.455 ;
        RECT  2.155 0.570 2.430 2.760 ;
        RECT  1.670 0.520 1.915 1.330 ;
        RECT  0.470 1.090 1.670 1.330 ;
        RECT  0.230 0.520 0.470 1.330 ;
    END
END CKLNQD1BWP7T

MACRO CKLNQD2BWP7T
    CLASS CORE ;
    FOREIGN CKLNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 1.0328 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.690 1.210 9.940 2.710 ;
        RECT  9.685 0.795 9.690 2.710 ;
        RECT  9.660 0.795 9.685 3.220 ;
        RECT  9.445 0.795 9.660 1.465 ;
        RECT  9.445 2.195 9.660 3.220 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.680 1.555 2.710 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.5859 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.660 7.140 2.710 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.415 -0.235 10.640 0.235 ;
        RECT  10.170 -0.235 10.415 1.165 ;
        RECT  8.965 -0.235 10.170 0.235 ;
        RECT  8.725 -0.235 8.965 1.190 ;
        RECT  5.515 -0.235 8.725 0.235 ;
        RECT  5.175 -0.235 5.515 0.465 ;
        RECT  3.885 -0.235 5.175 0.235 ;
        RECT  3.655 -0.235 3.885 0.860 ;
        RECT  1.265 -0.235 3.655 0.235 ;
        RECT  0.885 -0.235 1.265 0.820 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.410 3.685 10.640 4.155 ;
        RECT  10.175 2.245 10.410 4.155 ;
        RECT  9.030 3.685 10.175 4.155 ;
        RECT  8.650 3.030 9.030 4.155 ;
        RECT  7.315 3.685 8.650 4.155 ;
        RECT  6.975 3.245 7.315 4.155 ;
        RECT  5.895 3.685 6.975 4.155 ;
        RECT  5.515 2.870 5.895 4.155 ;
        RECT  3.615 3.685 5.515 4.155 ;
        RECT  3.380 2.995 3.615 4.155 ;
        RECT  0.540 3.685 3.380 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.930 1.600 9.160 2.530 ;
        RECT  8.245 2.290 8.930 2.530 ;
        RECT  8.245 0.465 8.485 1.970 ;
        RECT  6.055 0.465 8.245 0.705 ;
        RECT  8.005 2.290 8.245 3.335 ;
        RECT  7.890 2.290 8.005 2.530 ;
        RECT  7.660 0.935 7.890 2.530 ;
        RECT  7.130 0.935 7.660 1.175 ;
        RECT  6.595 0.935 6.715 1.180 ;
        RECT  6.365 0.935 6.595 3.050 ;
        RECT  6.315 2.030 6.365 3.050 ;
        RECT  5.315 2.030 6.315 2.270 ;
        RECT  5.815 0.465 6.055 0.925 ;
        RECT  4.610 0.695 5.815 0.925 ;
        RECT  5.085 1.170 5.375 1.420 ;
        RECT  4.830 1.170 5.085 3.455 ;
        RECT  4.075 3.225 4.830 3.455 ;
        RECT  4.600 0.515 4.610 0.925 ;
        RECT  4.370 0.515 4.600 2.760 ;
        RECT  4.310 1.995 4.370 2.760 ;
        RECT  3.425 1.995 4.310 2.225 ;
        RECT  3.425 1.235 4.125 1.575 ;
        RECT  3.845 2.495 4.075 3.455 ;
        RECT  2.965 2.495 3.845 2.725 ;
        RECT  3.195 0.570 3.425 1.575 ;
        RECT  3.195 1.855 3.425 2.225 ;
        RECT  2.430 0.570 3.195 0.805 ;
        RECT  2.735 1.115 2.965 3.455 ;
        RECT  1.850 3.215 2.735 3.455 ;
        RECT  2.155 0.570 2.430 2.760 ;
        RECT  1.670 0.520 1.915 1.330 ;
        RECT  0.470 1.090 1.670 1.330 ;
        RECT  0.230 0.520 0.470 1.330 ;
    END
END CKLNQD2BWP7T

MACRO CKLNQD4BWP7T
    CLASS CORE ;
    FOREIGN CKLNQD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 2.0466 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.240 0.490 12.490 3.205 ;
        RECT  11.590 0.990 12.240 2.550 ;
        RECT  11.055 0.990 11.590 1.340 ;
        RECT  11.055 2.200 11.590 2.550 ;
        RECT  10.805 0.490 11.055 1.340 ;
        RECT  10.800 2.200 11.055 3.205 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.680 1.555 2.710 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 0.8019 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.520 1.695 9.860 2.660 ;
        RECT  7.730 2.380 9.520 2.660 ;
        RECT  7.500 1.680 7.730 2.660 ;
        RECT  6.825 1.680 7.500 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.290 -0.235 13.440 0.235 ;
        RECT  12.910 -0.235 13.290 0.735 ;
        RECT  11.850 -0.235 12.910 0.235 ;
        RECT  11.470 -0.235 11.850 0.730 ;
        RECT  10.355 -0.235 11.470 0.235 ;
        RECT  9.975 -0.235 10.355 0.730 ;
        RECT  5.665 -0.235 9.975 0.235 ;
        RECT  5.325 -0.235 5.665 0.465 ;
        RECT  3.885 -0.235 5.325 0.235 ;
        RECT  3.655 -0.235 3.885 0.860 ;
        RECT  1.265 -0.235 3.655 0.235 ;
        RECT  0.885 -0.235 1.265 0.820 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.280 3.685 13.440 4.155 ;
        RECT  12.900 2.305 13.280 4.155 ;
        RECT  11.850 3.685 12.900 4.155 ;
        RECT  11.470 2.780 11.850 4.155 ;
        RECT  10.340 3.685 11.470 4.155 ;
        RECT  10.000 3.450 10.340 4.155 ;
        RECT  8.800 3.685 10.000 4.155 ;
        RECT  8.460 3.450 8.800 4.155 ;
        RECT  7.270 3.685 8.460 4.155 ;
        RECT  7.030 2.555 7.270 4.155 ;
        RECT  5.895 3.685 7.030 4.155 ;
        RECT  5.515 2.870 5.895 4.155 ;
        RECT  3.615 3.685 5.515 4.155 ;
        RECT  3.380 2.995 3.615 4.155 ;
        RECT  0.540 3.685 3.380 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.055 0.990 11.390 1.340 ;
        RECT  11.055 2.200 11.390 2.550 ;
        RECT  10.805 0.490 11.055 1.340 ;
        RECT  10.800 2.200 11.055 3.205 ;
        RECT  10.380 1.610 11.330 1.850 ;
        RECT  10.140 1.215 10.380 3.120 ;
        RECT  8.800 1.215 10.140 1.445 ;
        RECT  7.700 2.890 10.140 3.120 ;
        RECT  9.220 0.465 9.560 0.985 ;
        RECT  8.040 0.465 9.220 0.695 ;
        RECT  8.190 1.685 9.030 1.930 ;
        RECT  8.460 0.925 8.800 1.445 ;
        RECT  7.960 1.215 8.190 1.930 ;
        RECT  7.700 0.465 8.040 0.985 ;
        RECT  7.285 1.215 7.960 1.450 ;
        RECT  7.055 0.465 7.285 1.450 ;
        RECT  6.135 0.465 7.055 0.695 ;
        RECT  6.595 0.925 6.715 1.155 ;
        RECT  6.365 0.925 6.595 3.050 ;
        RECT  6.315 2.030 6.365 3.050 ;
        RECT  5.315 2.030 6.315 2.270 ;
        RECT  5.895 0.465 6.135 0.925 ;
        RECT  4.610 0.695 5.895 0.925 ;
        RECT  5.085 1.170 5.375 1.420 ;
        RECT  4.830 1.170 5.085 3.455 ;
        RECT  4.075 3.225 4.830 3.455 ;
        RECT  4.600 0.515 4.610 0.925 ;
        RECT  4.370 0.515 4.600 2.760 ;
        RECT  4.310 1.995 4.370 2.760 ;
        RECT  3.425 1.995 4.310 2.225 ;
        RECT  3.425 1.235 4.125 1.575 ;
        RECT  3.845 2.495 4.075 3.455 ;
        RECT  2.965 2.495 3.845 2.725 ;
        RECT  3.195 0.570 3.425 1.575 ;
        RECT  3.195 1.855 3.425 2.225 ;
        RECT  2.430 0.570 3.195 0.805 ;
        RECT  2.735 1.115 2.965 3.455 ;
        RECT  1.850 3.215 2.735 3.455 ;
        RECT  2.155 0.570 2.430 2.760 ;
        RECT  1.670 0.520 1.915 1.330 ;
        RECT  0.470 1.090 1.670 1.330 ;
        RECT  0.230 0.520 0.470 1.330 ;
    END
END CKLNQD4BWP7T

MACRO CKLNQD6BWP7T
    CLASS CORE ;
    FOREIGN CKLNQD6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 3.0699 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.055 0.640 15.290 1.405 ;
        RECT  15.055 2.155 15.290 3.200 ;
        RECT  14.730 1.175 15.055 1.405 ;
        RECT  14.730 2.155 15.055 2.505 ;
        RECT  13.850 1.175 14.730 2.505 ;
        RECT  13.830 0.640 13.850 3.200 ;
        RECT  13.615 0.640 13.830 1.405 ;
        RECT  13.615 2.155 13.830 3.200 ;
        RECT  12.410 1.175 13.615 1.405 ;
        RECT  12.410 2.155 13.615 2.505 ;
        RECT  12.170 0.660 12.410 1.405 ;
        RECT  12.175 2.155 12.410 3.200 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.680 1.555 2.710 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 1.0989 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.190 1.845 9.025 2.100 ;
        RECT  6.185 1.820 7.190 2.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.010 ;
        RECT  14.640 -0.235 15.775 0.235 ;
        RECT  14.260 -0.235 14.640 0.945 ;
        RECT  13.200 -0.235 14.260 0.235 ;
        RECT  12.820 -0.235 13.200 0.945 ;
        RECT  11.765 -0.235 12.820 0.235 ;
        RECT  11.385 -0.235 11.765 1.015 ;
        RECT  5.665 -0.235 11.385 0.235 ;
        RECT  5.325 -0.235 5.665 0.465 ;
        RECT  3.885 -0.235 5.325 0.235 ;
        RECT  3.655 -0.235 3.885 0.860 ;
        RECT  1.265 -0.235 3.655 0.235 ;
        RECT  0.885 -0.235 1.265 0.820 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.080 3.685 16.240 4.155 ;
        RECT  15.700 2.305 16.080 4.155 ;
        RECT  14.640 3.685 15.700 4.155 ;
        RECT  14.260 2.780 14.640 4.155 ;
        RECT  13.200 3.685 14.260 4.155 ;
        RECT  12.820 2.780 13.200 4.155 ;
        RECT  11.765 3.685 12.820 4.155 ;
        RECT  11.385 3.140 11.765 4.155 ;
        RECT  10.325 3.685 11.385 4.155 ;
        RECT  9.945 3.140 10.325 4.155 ;
        RECT  8.885 3.685 9.945 4.155 ;
        RECT  8.505 3.140 8.885 4.155 ;
        RECT  7.365 3.685 8.505 4.155 ;
        RECT  7.135 2.650 7.365 4.155 ;
        RECT  5.895 3.685 7.135 4.155 ;
        RECT  5.515 2.975 5.895 4.155 ;
        RECT  3.615 3.685 5.515 4.155 ;
        RECT  3.380 2.995 3.615 4.155 ;
        RECT  0.540 3.685 3.380 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.055 0.640 15.290 1.405 ;
        RECT  15.055 2.155 15.290 3.200 ;
        RECT  14.930 1.175 15.055 1.405 ;
        RECT  14.930 2.155 15.055 2.505 ;
        RECT  13.615 0.640 13.630 1.405 ;
        RECT  13.615 2.155 13.630 3.200 ;
        RECT  12.410 1.175 13.615 1.405 ;
        RECT  12.410 2.155 13.615 2.505 ;
        RECT  12.170 0.660 12.410 1.405 ;
        RECT  12.175 2.155 12.410 3.200 ;
        RECT  11.815 1.660 13.580 1.895 ;
        RECT  11.585 1.265 11.815 2.800 ;
        RECT  10.400 1.265 11.585 1.495 ;
        RECT  10.965 2.570 11.585 2.800 ;
        RECT  9.895 1.725 11.240 1.955 ;
        RECT  10.680 0.465 11.020 1.035 ;
        RECT  10.735 2.570 10.965 3.385 ;
        RECT  9.525 2.570 10.735 2.800 ;
        RECT  8.140 0.465 10.680 0.695 ;
        RECT  10.170 0.925 10.400 1.495 ;
        RECT  8.510 0.925 10.170 1.155 ;
        RECT  9.665 1.385 9.895 1.955 ;
        RECT  7.570 1.385 9.665 1.615 ;
        RECT  9.295 2.570 9.525 3.385 ;
        RECT  8.085 2.570 9.295 2.800 ;
        RECT  7.800 0.465 8.140 1.035 ;
        RECT  7.800 2.570 8.085 3.385 ;
        RECT  7.340 0.465 7.570 1.615 ;
        RECT  6.135 0.465 7.340 0.695 ;
        RECT  6.430 0.965 6.660 1.485 ;
        RECT  6.330 2.515 6.560 3.195 ;
        RECT  5.895 1.255 6.430 1.485 ;
        RECT  5.600 2.515 6.330 2.745 ;
        RECT  5.895 0.465 6.135 0.925 ;
        RECT  4.610 0.695 5.895 0.925 ;
        RECT  5.665 1.255 5.895 1.880 ;
        RECT  5.600 1.650 5.665 1.880 ;
        RECT  5.370 1.650 5.600 2.745 ;
        RECT  5.085 1.170 5.375 1.420 ;
        RECT  4.830 1.170 5.085 3.455 ;
        RECT  4.075 3.225 4.830 3.455 ;
        RECT  4.600 0.515 4.610 0.925 ;
        RECT  4.370 0.515 4.600 2.760 ;
        RECT  4.310 1.995 4.370 2.760 ;
        RECT  3.425 1.995 4.310 2.225 ;
        RECT  3.425 1.235 4.125 1.575 ;
        RECT  3.845 2.495 4.075 3.455 ;
        RECT  2.965 2.495 3.845 2.725 ;
        RECT  3.195 0.570 3.425 1.575 ;
        RECT  3.195 1.855 3.425 2.225 ;
        RECT  2.430 0.570 3.195 0.805 ;
        RECT  2.735 1.115 2.965 3.455 ;
        RECT  1.850 3.215 2.735 3.455 ;
        RECT  2.155 0.570 2.430 2.760 ;
        RECT  1.670 0.520 1.915 1.330 ;
        RECT  0.470 1.090 1.670 1.330 ;
        RECT  0.230 0.520 0.470 1.330 ;
    END
END CKLNQD6BWP7T

MACRO CKLNQD8BWP7T
    CLASS CORE ;
    FOREIGN CKLNQD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN TE
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END TE
    PIN Q
        ANTENNADIFFAREA 4.5639 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.335 0.485 16.570 1.160 ;
        RECT  16.330 2.180 16.570 3.135 ;
        RECT  15.290 0.905 16.335 1.160 ;
        RECT  15.290 2.180 16.330 2.530 ;
        RECT  15.130 0.905 15.290 2.530 ;
        RECT  14.895 0.595 15.130 3.135 ;
        RECT  14.890 0.905 14.895 3.135 ;
        RECT  14.390 0.905 14.890 2.530 ;
        RECT  13.690 0.905 14.390 1.160 ;
        RECT  13.690 2.180 14.390 2.530 ;
        RECT  13.455 0.595 13.690 1.160 ;
        RECT  13.450 2.180 13.690 3.135 ;
        RECT  12.250 0.905 13.455 1.160 ;
        RECT  12.250 2.180 13.450 2.530 ;
        RECT  12.010 0.490 12.250 1.160 ;
        RECT  12.010 2.180 12.250 3.135 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.680 1.555 2.710 ;
        END
    END E
    PIN CP
        ANTENNAGATEAREA 1.1097 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.260 1.845 8.920 2.100 ;
        RECT  6.220 1.820 7.260 2.100 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.920 -0.235 16.800 0.235 ;
        RECT  15.540 -0.235 15.920 0.675 ;
        RECT  14.480 -0.235 15.540 0.235 ;
        RECT  14.100 -0.235 14.480 0.675 ;
        RECT  13.040 -0.235 14.100 0.235 ;
        RECT  12.660 -0.235 13.040 0.675 ;
        RECT  11.600 -0.235 12.660 0.235 ;
        RECT  11.220 -0.235 11.600 0.670 ;
        RECT  5.665 -0.235 11.220 0.235 ;
        RECT  5.325 -0.235 5.665 0.465 ;
        RECT  3.885 -0.235 5.325 0.235 ;
        RECT  3.655 -0.235 3.885 0.860 ;
        RECT  1.265 -0.235 3.655 0.235 ;
        RECT  0.885 -0.235 1.265 0.820 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.920 3.685 16.800 4.155 ;
        RECT  15.540 2.775 15.920 4.155 ;
        RECT  14.480 3.685 15.540 4.155 ;
        RECT  14.100 2.775 14.480 4.155 ;
        RECT  13.040 3.685 14.100 4.155 ;
        RECT  12.660 2.775 13.040 4.155 ;
        RECT  11.600 3.685 12.660 4.155 ;
        RECT  11.220 3.140 11.600 4.155 ;
        RECT  10.160 3.685 11.220 4.155 ;
        RECT  9.780 3.140 10.160 4.155 ;
        RECT  8.720 3.685 9.780 4.155 ;
        RECT  8.340 3.140 8.720 4.155 ;
        RECT  7.280 3.685 8.340 4.155 ;
        RECT  6.900 3.210 7.280 4.155 ;
        RECT  5.895 3.685 6.900 4.155 ;
        RECT  5.515 2.860 5.895 4.155 ;
        RECT  3.615 3.685 5.515 4.155 ;
        RECT  3.380 2.995 3.615 4.155 ;
        RECT  0.540 3.685 3.380 4.155 ;
        RECT  0.160 3.040 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.335 0.485 16.570 1.160 ;
        RECT  16.330 2.180 16.570 3.135 ;
        RECT  15.490 0.905 16.335 1.160 ;
        RECT  15.490 2.180 16.330 2.530 ;
        RECT  13.690 0.905 14.190 1.160 ;
        RECT  13.690 2.180 14.190 2.530 ;
        RECT  13.455 0.595 13.690 1.160 ;
        RECT  13.450 2.180 13.690 3.135 ;
        RECT  12.250 0.905 13.455 1.160 ;
        RECT  12.250 2.180 13.450 2.530 ;
        RECT  12.010 0.490 12.250 1.160 ;
        RECT  12.010 2.180 12.250 3.135 ;
        RECT  11.650 1.450 13.885 1.695 ;
        RECT  11.420 1.295 11.650 2.800 ;
        RECT  10.235 1.295 11.420 1.525 ;
        RECT  10.800 2.570 11.420 2.800 ;
        RECT  9.730 1.755 11.075 1.985 ;
        RECT  10.475 0.465 10.815 1.065 ;
        RECT  10.570 2.570 10.800 3.385 ;
        RECT  9.360 2.570 10.570 2.800 ;
        RECT  7.975 0.465 10.475 0.695 ;
        RECT  10.005 0.925 10.235 1.525 ;
        RECT  8.305 0.925 10.005 1.155 ;
        RECT  9.500 1.385 9.730 1.985 ;
        RECT  8.105 1.385 9.500 1.615 ;
        RECT  9.130 2.570 9.360 3.385 ;
        RECT  7.920 2.570 9.130 2.800 ;
        RECT  7.875 1.295 8.105 1.615 ;
        RECT  7.635 0.465 7.975 1.065 ;
        RECT  7.635 2.570 7.920 3.385 ;
        RECT  7.275 1.295 7.875 1.525 ;
        RECT  7.045 0.465 7.275 1.525 ;
        RECT  6.135 0.465 7.045 0.695 ;
        RECT  6.430 0.955 6.660 1.385 ;
        RECT  6.315 2.400 6.595 2.880 ;
        RECT  5.935 1.155 6.430 1.385 ;
        RECT  5.600 2.400 6.315 2.630 ;
        RECT  5.895 0.465 6.135 0.925 ;
        RECT  5.705 1.155 5.935 1.880 ;
        RECT  4.610 0.695 5.895 0.925 ;
        RECT  5.600 1.650 5.705 1.880 ;
        RECT  5.370 1.650 5.600 2.630 ;
        RECT  5.085 1.170 5.375 1.420 ;
        RECT  4.830 1.170 5.085 3.455 ;
        RECT  4.075 3.225 4.830 3.455 ;
        RECT  4.600 0.515 4.610 0.925 ;
        RECT  4.370 0.515 4.600 2.760 ;
        RECT  4.310 1.995 4.370 2.760 ;
        RECT  3.425 1.995 4.310 2.225 ;
        RECT  3.425 1.235 4.125 1.575 ;
        RECT  3.845 2.495 4.075 3.455 ;
        RECT  2.965 2.495 3.845 2.725 ;
        RECT  3.195 0.570 3.425 1.575 ;
        RECT  3.195 1.855 3.425 2.225 ;
        RECT  2.430 0.570 3.195 0.805 ;
        RECT  2.735 1.115 2.965 3.455 ;
        RECT  1.850 3.215 2.735 3.455 ;
        RECT  2.155 0.570 2.430 2.760 ;
        RECT  1.670 0.520 1.915 1.330 ;
        RECT  0.470 1.090 1.670 1.330 ;
        RECT  0.230 0.520 0.470 1.330 ;
    END
END CKLNQD8BWP7T

MACRO CKMUX2D0BWP7T
    CLASS CORE ;
    FOREIGN CKMUX2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.6432 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 0.465 4.900 3.220 ;
        RECT  4.520 0.465 4.620 0.695 ;
        RECT  4.570 2.365 4.620 3.220 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.5751 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 0.930 3.045 1.270 ;
        RECT  2.720 0.930 2.950 1.695 ;
        RECT  2.425 1.465 2.720 1.695 ;
        RECT  2.195 1.465 2.425 2.455 ;
        RECT  1.990 2.225 2.195 2.455 ;
        RECT  1.760 2.225 1.990 2.610 ;
        RECT  0.980 2.380 1.760 2.610 ;
        RECT  0.700 1.210 0.980 2.610 ;
        RECT  0.575 1.570 0.700 2.040 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.2961 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 1.210 3.780 2.190 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2961 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.210 1.540 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.120 -0.235 5.040 0.235 ;
        RECT  3.740 -0.235 4.120 0.510 ;
        RECT  1.280 -0.235 3.740 0.235 ;
        RECT  0.940 -0.235 1.280 0.465 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 3.685 5.040 4.155 ;
        RECT  3.800 2.945 4.140 4.155 ;
        RECT  1.285 3.685 3.800 4.155 ;
        RECT  0.945 3.320 1.285 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.295 1.640 4.385 1.980 ;
        RECT  4.065 0.745 4.295 2.715 ;
        RECT  3.510 0.745 4.065 0.980 ;
        RECT  3.485 2.485 4.065 2.715 ;
        RECT  3.275 0.465 3.510 0.980 ;
        RECT  3.255 2.485 3.485 3.455 ;
        RECT  2.380 0.465 3.275 0.695 ;
        RECT  2.650 3.225 3.255 3.455 ;
        RECT  3.025 1.925 3.230 2.155 ;
        RECT  2.795 1.925 3.025 2.995 ;
        RECT  2.410 2.765 2.795 2.995 ;
        RECT  2.155 0.985 2.430 1.215 ;
        RECT  2.180 2.765 2.410 3.070 ;
        RECT  0.345 2.840 2.180 3.070 ;
        RECT  1.925 0.750 2.155 1.215 ;
        RECT  0.520 0.750 1.925 0.980 ;
        RECT  0.345 0.465 0.520 0.980 ;
        RECT  0.115 0.465 0.345 3.070 ;
    END
END CKMUX2D0BWP7T

MACRO CKMUX2D1BWP7T
    CLASS CORE ;
    FOREIGN CKMUX2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.9936 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 0.465 4.900 3.220 ;
        RECT  4.520 0.465 4.620 0.695 ;
        RECT  4.570 2.365 4.620 3.220 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.6714 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.690 1.000 2.905 1.340 ;
        RECT  2.460 1.000 2.690 1.745 ;
        RECT  2.425 1.515 2.460 1.745 ;
        RECT  2.195 1.515 2.425 2.455 ;
        RECT  1.990 2.225 2.195 2.455 ;
        RECT  1.760 2.225 1.990 2.610 ;
        RECT  0.980 2.380 1.760 2.610 ;
        RECT  0.700 1.210 0.980 2.610 ;
        RECT  0.575 1.570 0.700 2.040 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.3303 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 1.155 3.780 2.190 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3303 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.210 1.540 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.120 -0.235 5.040 0.235 ;
        RECT  3.740 -0.235 4.120 0.465 ;
        RECT  1.280 -0.235 3.740 0.235 ;
        RECT  0.940 -0.235 1.280 0.465 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 3.685 5.040 4.155 ;
        RECT  3.800 3.155 4.140 4.155 ;
        RECT  1.280 3.685 3.800 4.155 ;
        RECT  0.940 3.450 1.280 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.290 1.725 4.385 2.065 ;
        RECT  4.060 0.695 4.290 2.925 ;
        RECT  3.510 0.695 4.060 0.925 ;
        RECT  3.485 2.695 4.060 2.925 ;
        RECT  3.275 0.465 3.510 0.925 ;
        RECT  3.255 2.695 3.485 3.455 ;
        RECT  2.380 0.465 3.275 0.695 ;
        RECT  2.630 3.225 3.255 3.455 ;
        RECT  3.025 1.725 3.155 2.280 ;
        RECT  2.925 1.725 3.025 2.995 ;
        RECT  2.795 2.050 2.925 2.995 ;
        RECT  2.390 2.765 2.795 2.995 ;
        RECT  2.160 2.765 2.390 3.170 ;
        RECT  2.010 1.055 2.230 1.285 ;
        RECT  0.470 2.940 2.160 3.170 ;
        RECT  1.780 0.750 2.010 1.285 ;
        RECT  0.520 0.750 1.780 0.980 ;
        RECT  0.345 0.465 0.520 0.980 ;
        RECT  0.345 2.795 0.470 3.170 ;
        RECT  0.115 0.465 0.345 3.170 ;
    END
END CKMUX2D1BWP7T

MACRO CKMUX2D2BWP7T
    CLASS CORE ;
    FOREIGN CKMUX2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1322 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 0.495 5.460 2.600 ;
        RECT  5.180 0.495 5.205 3.370 ;
        RECT  4.975 0.495 5.180 0.835 ;
        RECT  4.975 2.350 5.180 3.370 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.7605 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.595 1.385 2.825 1.905 ;
        RECT  2.560 1.675 2.595 1.905 ;
        RECT  2.330 1.675 2.560 3.020 ;
        RECT  0.980 2.790 2.330 3.020 ;
        RECT  0.700 1.445 0.980 3.020 ;
        RECT  0.575 1.445 0.700 2.035 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4194 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.005 1.375 4.240 2.000 ;
        RECT  3.780 1.770 4.005 2.000 ;
        RECT  3.500 1.770 3.780 2.710 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.4194 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.770 2.100 2.150 ;
        RECT  1.250 1.385 1.540 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 -0.235 6.160 0.235 ;
        RECT  5.695 -0.235 5.925 0.935 ;
        RECT  4.500 -0.235 5.695 0.235 ;
        RECT  4.160 -0.235 4.500 0.465 ;
        RECT  1.280 -0.235 4.160 0.235 ;
        RECT  0.940 -0.235 1.280 0.675 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 3.685 6.160 4.155 ;
        RECT  5.695 2.245 5.925 4.155 ;
        RECT  4.500 3.685 5.695 4.155 ;
        RECT  4.160 3.455 4.500 4.155 ;
        RECT  1.280 3.685 4.160 4.155 ;
        RECT  0.900 3.250 1.280 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.745 1.375 4.940 1.715 ;
        RECT  4.515 0.695 4.745 3.225 ;
        RECT  3.930 0.695 4.515 0.925 ;
        RECT  3.180 2.995 4.515 3.225 ;
        RECT  3.695 0.465 3.930 0.925 ;
        RECT  2.275 0.465 3.695 0.695 ;
        RECT  3.285 1.110 3.495 1.450 ;
        RECT  3.055 0.925 3.285 1.450 ;
        RECT  2.945 2.150 3.180 3.225 ;
        RECT  2.210 0.925 3.055 1.155 ;
        RECT  1.870 0.925 2.210 1.395 ;
        RECT  0.465 0.925 1.870 1.155 ;
        RECT  0.345 2.375 0.470 3.285 ;
        RECT  0.345 0.495 0.465 1.155 ;
        RECT  0.115 0.495 0.345 3.285 ;
    END
END CKMUX2D2BWP7T

MACRO CKND0BWP7T
    CLASS CORE ;
    FOREIGN CKND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.8215 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 0.545 1.540 3.405 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2790 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.605 0.915 1.945 ;
        RECT  0.140 1.605 0.420 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 -0.235 1.680 0.235 ;
        RECT  0.320 -0.235 0.700 0.925 ;
        RECT  0.000 -0.235 0.320 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 3.685 1.680 4.155 ;
        RECT  0.320 3.020 0.700 4.155 ;
        RECT  0.000 3.685 0.320 4.155 ;
        END
    END VDD
END CKND0BWP7T

MACRO CKND10BWP7T
    CLASS CORE ;
    FOREIGN CKND10BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.4158 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.705 2.105 6.960 3.380 ;
        RECT  5.520 2.105 6.705 2.505 ;
        RECT  5.990 0.505 6.230 1.310 ;
        RECT  4.790 0.910 5.990 1.310 ;
        RECT  5.265 2.105 5.520 3.310 ;
        RECT  4.650 2.105 5.265 2.505 ;
        RECT  4.650 0.505 4.790 1.310 ;
        RECT  4.550 0.505 4.650 2.505 ;
        RECT  4.080 0.910 4.550 2.505 ;
        RECT  3.825 0.910 4.080 3.310 ;
        RECT  3.350 0.910 3.825 2.505 ;
        RECT  3.190 0.505 3.350 2.505 ;
        RECT  3.110 0.505 3.190 1.310 ;
        RECT  2.640 2.105 3.190 2.505 ;
        RECT  1.910 0.910 3.110 1.310 ;
        RECT  2.385 2.105 2.640 3.310 ;
        RECT  1.200 2.105 2.385 2.505 ;
        RECT  1.670 0.505 1.910 1.310 ;
        RECT  0.945 2.105 1.200 3.380 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 3.4083 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.540 2.890 1.770 ;
        RECT  0.140 0.620 0.465 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.020 -0.235 7.280 0.235 ;
        RECT  6.640 -0.235 7.020 0.810 ;
        RECT  5.630 -0.235 6.640 0.235 ;
        RECT  5.170 -0.235 5.630 0.670 ;
        RECT  4.190 -0.235 5.170 0.235 ;
        RECT  3.730 -0.235 4.190 0.670 ;
        RECT  2.750 -0.235 3.730 0.235 ;
        RECT  2.290 -0.235 2.750 0.670 ;
        RECT  1.270 -0.235 2.290 0.235 ;
        RECT  0.890 -0.235 1.270 0.800 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.310 3.685 7.280 4.155 ;
        RECT  5.925 2.780 6.310 4.155 ;
        RECT  4.870 3.685 5.925 4.155 ;
        RECT  4.485 2.780 4.870 4.155 ;
        RECT  3.430 3.685 4.485 4.155 ;
        RECT  3.045 2.780 3.430 4.155 ;
        RECT  1.990 3.685 3.045 4.155 ;
        RECT  1.605 2.780 1.990 4.155 ;
        RECT  0.540 3.685 1.605 4.155 ;
        RECT  0.160 2.570 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.705 2.105 6.960 3.380 ;
        RECT  5.520 2.105 6.705 2.505 ;
        RECT  5.990 0.505 6.230 1.310 ;
        RECT  4.850 0.910 5.990 1.310 ;
        RECT  5.265 2.105 5.520 3.310 ;
        RECT  4.850 2.105 5.265 2.505 ;
        RECT  1.910 0.910 2.990 1.310 ;
        RECT  2.640 2.105 2.990 2.505 ;
        RECT  2.385 2.105 2.640 3.310 ;
        RECT  1.200 2.105 2.385 2.505 ;
        RECT  1.670 0.505 1.910 1.310 ;
        RECT  0.945 2.105 1.200 3.380 ;
    END
END CKND10BWP7T

MACRO CKND12BWP7T
    CLASS CORE ;
    FOREIGN CKND12BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 6.4300 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.145 2.105 8.400 3.375 ;
        RECT  6.960 2.105 8.145 2.505 ;
        RECT  7.430 0.610 7.670 1.375 ;
        RECT  6.230 0.975 7.430 1.375 ;
        RECT  6.705 2.105 6.960 3.365 ;
        RECT  5.520 2.105 6.705 2.505 ;
        RECT  5.990 0.610 6.230 1.375 ;
        RECT  5.210 0.975 5.990 1.375 ;
        RECT  5.265 2.105 5.520 3.365 ;
        RECT  5.210 2.105 5.265 2.505 ;
        RECT  4.790 0.975 5.210 2.505 ;
        RECT  4.550 0.610 4.790 2.505 ;
        RECT  4.080 0.975 4.550 2.505 ;
        RECT  3.825 0.975 4.080 3.365 ;
        RECT  3.750 0.975 3.825 2.505 ;
        RECT  3.350 0.975 3.750 1.375 ;
        RECT  2.640 2.105 3.750 2.505 ;
        RECT  3.110 0.610 3.350 1.375 ;
        RECT  1.910 0.975 3.110 1.375 ;
        RECT  2.385 2.105 2.640 3.365 ;
        RECT  1.200 2.105 2.385 2.505 ;
        RECT  1.670 0.570 1.910 1.375 ;
        RECT  0.945 2.105 1.200 3.365 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 4.0932 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.615 3.360 1.875 ;
        RECT  0.140 0.750 0.465 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.460 -0.235 8.960 0.235 ;
        RECT  8.080 -0.235 8.460 0.840 ;
        RECT  7.020 -0.235 8.080 0.235 ;
        RECT  6.640 -0.235 7.020 0.735 ;
        RECT  5.590 -0.235 6.640 0.235 ;
        RECT  5.210 -0.235 5.590 0.735 ;
        RECT  4.150 -0.235 5.210 0.235 ;
        RECT  3.770 -0.235 4.150 0.735 ;
        RECT  2.710 -0.235 3.770 0.235 ;
        RECT  2.330 -0.235 2.710 0.735 ;
        RECT  1.270 -0.235 2.330 0.235 ;
        RECT  0.890 -0.235 1.270 0.840 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.750 3.685 8.960 4.155 ;
        RECT  7.365 2.780 7.750 4.155 ;
        RECT  6.310 3.685 7.365 4.155 ;
        RECT  5.925 2.780 6.310 4.155 ;
        RECT  4.870 3.685 5.925 4.155 ;
        RECT  4.485 2.780 4.870 4.155 ;
        RECT  3.430 3.685 4.485 4.155 ;
        RECT  3.045 2.780 3.430 4.155 ;
        RECT  1.990 3.685 3.045 4.155 ;
        RECT  1.605 2.780 1.990 4.155 ;
        RECT  0.540 3.685 1.605 4.155 ;
        RECT  0.160 2.520 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.145 2.105 8.400 3.375 ;
        RECT  6.960 2.105 8.145 2.505 ;
        RECT  7.430 0.610 7.670 1.375 ;
        RECT  6.230 0.975 7.430 1.375 ;
        RECT  6.705 2.105 6.960 3.365 ;
        RECT  5.520 2.105 6.705 2.505 ;
        RECT  5.990 0.610 6.230 1.375 ;
        RECT  5.410 0.975 5.990 1.375 ;
        RECT  5.410 2.105 5.520 3.365 ;
        RECT  3.350 0.975 3.550 1.375 ;
        RECT  2.640 2.105 3.550 2.505 ;
        RECT  3.110 0.610 3.350 1.375 ;
        RECT  1.910 0.975 3.110 1.375 ;
        RECT  2.385 2.105 2.640 3.365 ;
        RECT  1.200 2.105 2.385 2.505 ;
        RECT  1.670 0.570 1.910 1.375 ;
        RECT  0.945 2.105 1.200 3.365 ;
    END
END CKND12BWP7T

MACRO CKND1BWP7T
    CLASS CORE ;
    FOREIGN CKND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.0044 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 0.530 1.540 3.390 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.3411 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.605 0.915 1.945 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 -0.235 1.680 0.235 ;
        RECT  0.320 -0.235 0.700 0.825 ;
        RECT  0.000 -0.235 0.320 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 3.685 1.680 4.155 ;
        RECT  0.320 2.455 0.700 4.155 ;
        RECT  0.000 3.685 0.320 4.155 ;
        END
    END VDD
END CKND1BWP7T

MACRO CKND2BWP7T
    CLASS CORE ;
    FOREIGN CKND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.0233 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.710 ;
        RECT  1.235 1.210 1.260 1.440 ;
        RECT  1.235 2.370 1.260 2.710 ;
        RECT  1.005 0.540 1.235 1.440 ;
        RECT  1.005 2.370 1.235 3.435 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.6822 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.660 0.935 1.890 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.080 0.830 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.815 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 3.685 2.240 4.155 ;
        RECT  1.775 2.245 2.005 4.155 ;
        RECT  0.540 3.685 1.775 4.155 ;
        RECT  0.160 2.500 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
END CKND2BWP7T

MACRO CKND2D0BWP7T
    CLASS CORE ;
    FOREIGN CKND2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6808 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.715 2.100 2.680 ;
        RECT  1.600 0.715 1.820 0.955 ;
        RECT  1.235 2.430 1.820 2.680 ;
        RECT  0.995 2.430 1.235 3.350 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2196 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.655 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2304 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.240 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.590 -0.235 2.240 0.235 ;
        RECT  0.210 -0.235 0.590 0.905 ;
        RECT  0.000 -0.235 0.210 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 3.685 2.240 4.155 ;
        RECT  1.655 3.080 2.035 4.155 ;
        RECT  0.590 3.685 1.655 4.155 ;
        RECT  0.210 3.080 0.590 4.155 ;
        RECT  0.000 3.685 0.210 4.155 ;
        END
    END VDD
END CKND2D0BWP7T

MACRO CKND2D1BWP7T
    CLASS CORE ;
    FOREIGN CKND2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2667 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.665 2.100 2.710 ;
        RECT  1.680 0.665 1.820 0.905 ;
        RECT  1.235 2.460 1.820 2.710 ;
        RECT  0.995 2.460 1.235 3.370 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.3699 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.655 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.240 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.590 -0.235 2.240 0.235 ;
        RECT  0.210 -0.235 0.590 0.830 ;
        RECT  0.000 -0.235 0.210 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 3.685 2.240 4.155 ;
        RECT  1.655 2.970 2.035 4.155 ;
        RECT  0.590 3.685 1.655 4.155 ;
        RECT  0.210 2.575 0.590 4.155 ;
        RECT  0.000 3.685 0.210 4.155 ;
        END
    END VDD
END CKND2D1BWP7T

MACRO CKND2D2BWP7T
    CLASS CORE ;
    FOREIGN CKND2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.0852 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.935 3.220 2.710 ;
        RECT  2.940 0.935 2.970 3.370 ;
        RECT  2.680 0.935 2.940 1.175 ;
        RECT  2.730 2.380 2.940 3.370 ;
        RECT  1.230 2.380 2.730 2.710 ;
        RECT  0.990 2.380 1.230 3.370 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.7092 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.655 1.520 1.900 ;
        RECT  0.140 1.655 0.420 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.7812 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.600 2.710 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 -0.235 3.920 0.235 ;
        RECT  0.920 -0.235 1.300 0.875 ;
        RECT  0.000 -0.235 0.920 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.690 3.685 3.920 4.155 ;
        RECT  3.450 2.250 3.690 4.155 ;
        RECT  2.130 3.685 3.450 4.155 ;
        RECT  1.750 2.950 2.130 4.155 ;
        RECT  0.590 3.685 1.750 4.155 ;
        RECT  0.210 2.950 0.590 4.155 ;
        RECT  0.000 3.685 0.210 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.450 0.465 3.690 1.305 ;
        RECT  2.060 0.465 3.450 0.705 ;
        RECT  1.820 0.465 2.060 1.335 ;
        RECT  0.510 1.105 1.820 1.335 ;
        RECT  0.270 0.760 0.510 1.335 ;
    END
END CKND2D2BWP7T

MACRO CKND2D3BWP7T
    CLASS CORE ;
    FOREIGN CKND2D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0514 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.570 0.575 4.815 1.380 ;
        RECT  4.090 1.040 4.570 1.380 ;
        RECT  3.830 1.040 4.090 3.120 ;
        RECT  3.405 1.040 3.830 2.750 ;
        RECT  3.190 0.925 3.405 2.750 ;
        RECT  3.065 0.925 3.190 1.380 ;
        RECT  2.630 2.400 3.190 2.750 ;
        RECT  2.390 2.400 2.630 3.240 ;
        RECT  1.190 2.400 2.390 2.750 ;
        RECT  0.950 2.400 1.190 3.240 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.0638 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.430 1.740 2.160 2.150 ;
        RECT  0.150 1.210 0.430 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.1718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.685 4.900 2.710 ;
        RECT  4.350 1.685 4.620 1.925 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.980 -0.235 5.040 0.235 ;
        RECT  1.600 -0.235 1.980 0.915 ;
        RECT  0.540 -0.235 1.600 0.235 ;
        RECT  0.160 -0.235 0.540 0.915 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.865 3.685 5.040 4.155 ;
        RECT  4.485 3.040 4.865 4.155 ;
        RECT  3.420 3.685 4.485 4.155 ;
        RECT  3.040 3.040 3.420 4.155 ;
        RECT  1.980 3.685 3.040 4.155 ;
        RECT  1.600 3.040 1.980 4.155 ;
        RECT  0.540 3.685 1.600 4.155 ;
        RECT  0.160 2.475 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.800 0.465 4.140 0.775 ;
        RECT  2.635 0.465 3.800 0.695 ;
        RECT  2.385 0.465 2.635 1.440 ;
        RECT  1.195 1.210 2.385 1.440 ;
        RECT  0.950 0.625 1.195 1.440 ;
    END
END CKND2D3BWP7T

MACRO CKND2D4BWP7T
    CLASS CORE ;
    FOREIGN CKND2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.8340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.325 0.925 5.665 1.455 ;
        RECT  5.375 2.430 5.615 3.240 ;
        RECT  4.650 2.430 5.375 2.780 ;
        RECT  4.650 1.225 5.325 1.455 ;
        RECT  4.225 1.225 4.650 2.780 ;
        RECT  4.180 0.925 4.225 2.780 ;
        RECT  3.930 0.925 4.180 3.240 ;
        RECT  3.885 0.925 3.930 2.780 ;
        RECT  3.750 1.225 3.885 2.780 ;
        RECT  2.735 2.430 3.750 2.780 ;
        RECT  2.485 2.430 2.735 3.240 ;
        RECT  1.295 2.430 2.485 2.780 ;
        RECT  1.045 2.430 1.295 3.240 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.4184 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.810 1.780 3.010 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.5624 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.025 1.695 6.070 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.800 -0.235 6.720 0.235 ;
        RECT  2.420 -0.235 2.800 0.780 ;
        RECT  1.360 -0.235 2.420 0.235 ;
        RECT  0.980 -0.235 1.360 0.780 ;
        RECT  0.000 -0.235 0.980 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.405 3.685 6.720 4.155 ;
        RECT  6.025 2.480 6.405 4.155 ;
        RECT  4.965 3.685 6.025 4.155 ;
        RECT  4.585 3.045 4.965 4.155 ;
        RECT  3.520 3.685 4.585 4.155 ;
        RECT  3.140 3.045 3.520 4.155 ;
        RECT  2.080 3.685 3.140 4.155 ;
        RECT  1.700 3.045 2.080 4.155 ;
        RECT  0.565 3.685 1.700 4.155 ;
        RECT  0.330 2.250 0.565 4.155 ;
        RECT  0.000 3.685 0.330 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.325 0.925 5.665 1.455 ;
        RECT  5.375 2.430 5.615 3.240 ;
        RECT  4.850 2.430 5.375 2.780 ;
        RECT  4.850 1.225 5.325 1.455 ;
        RECT  2.735 2.430 3.550 2.780 ;
        RECT  2.485 2.430 2.735 3.240 ;
        RECT  1.295 2.430 2.485 2.780 ;
        RECT  1.045 2.430 1.295 3.240 ;
        RECT  6.095 0.465 6.335 0.920 ;
        RECT  4.945 0.465 6.095 0.695 ;
        RECT  4.605 0.465 4.945 0.775 ;
        RECT  3.450 0.465 4.605 0.695 ;
        RECT  3.210 0.465 3.450 1.360 ;
        RECT  2.010 1.040 3.210 1.360 ;
        RECT  1.770 0.620 2.010 1.360 ;
        RECT  0.570 1.040 1.770 1.360 ;
        RECT  0.330 0.610 0.570 1.360 ;
    END
END CKND2D4BWP7T

MACRO CKND2D8BWP7T
    CLASS CORE ;
    FOREIGN CKND2D8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 8.0902 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.450 0.995 11.345 1.395 ;
        RECT  11.050 2.380 11.295 3.290 ;
        RECT  9.855 2.380 11.050 2.780 ;
        RECT  9.610 2.380 9.855 3.290 ;
        RECT  8.415 2.380 9.610 2.780 ;
        RECT  8.170 2.380 8.415 3.290 ;
        RECT  7.450 2.380 8.170 2.780 ;
        RECT  6.970 0.995 7.450 2.780 ;
        RECT  6.725 0.995 6.970 3.290 ;
        RECT  6.550 0.995 6.725 2.780 ;
        RECT  5.530 2.380 6.550 2.780 ;
        RECT  5.285 2.380 5.530 3.290 ;
        RECT  4.090 2.380 5.285 2.780 ;
        RECT  3.845 2.380 4.090 3.290 ;
        RECT  2.650 2.380 3.845 2.780 ;
        RECT  2.405 2.380 2.650 3.290 ;
        RECT  1.210 2.380 2.405 2.780 ;
        RECT  0.965 2.380 1.210 3.290 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 2.9520 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.740 5.790 1.970 ;
        RECT  0.700 1.740 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 3.4128 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.170 1.740 11.110 2.110 ;
        RECT  7.710 1.740 10.170 1.970 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.600 -0.235 12.320 0.235 ;
        RECT  5.220 -0.235 5.600 0.790 ;
        RECT  4.160 -0.235 5.220 0.235 ;
        RECT  3.780 -0.235 4.160 0.790 ;
        RECT  2.720 -0.235 3.780 0.235 ;
        RECT  2.340 -0.235 2.720 0.790 ;
        RECT  1.280 -0.235 2.340 0.235 ;
        RECT  0.900 -0.235 1.280 0.790 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.065 3.685 12.320 4.155 ;
        RECT  11.725 2.300 12.065 4.155 ;
        RECT  10.645 3.685 11.725 4.155 ;
        RECT  10.265 3.035 10.645 4.155 ;
        RECT  9.205 3.685 10.265 4.155 ;
        RECT  8.825 3.035 9.205 4.155 ;
        RECT  7.765 3.685 8.825 4.155 ;
        RECT  7.385 3.035 7.765 4.155 ;
        RECT  6.320 3.685 7.385 4.155 ;
        RECT  5.940 3.035 6.320 4.155 ;
        RECT  4.880 3.685 5.940 4.155 ;
        RECT  4.500 3.035 4.880 4.155 ;
        RECT  3.440 3.685 4.500 4.155 ;
        RECT  3.060 3.035 3.440 4.155 ;
        RECT  2.000 3.685 3.060 4.155 ;
        RECT  1.620 3.035 2.000 4.155 ;
        RECT  0.540 3.685 1.620 4.155 ;
        RECT  0.200 2.450 0.540 4.155 ;
        RECT  0.000 3.685 0.200 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.650 0.995 11.345 1.395 ;
        RECT  11.050 2.380 11.295 3.290 ;
        RECT  9.855 2.380 11.050 2.780 ;
        RECT  9.610 2.380 9.855 3.290 ;
        RECT  8.415 2.380 9.610 2.780 ;
        RECT  8.170 2.380 8.415 3.290 ;
        RECT  7.650 2.380 8.170 2.780 ;
        RECT  5.530 2.380 6.350 2.780 ;
        RECT  5.285 2.380 5.530 3.290 ;
        RECT  4.090 2.380 5.285 2.780 ;
        RECT  3.845 2.380 4.090 3.290 ;
        RECT  4.565 0.545 4.815 1.365 ;
        RECT  3.375 1.070 4.565 1.365 ;
        RECT  3.125 0.545 3.375 1.365 ;
        RECT  1.935 1.070 3.125 1.365 ;
        RECT  1.685 0.545 1.935 1.365 ;
        RECT  0.495 1.070 1.685 1.365 ;
        RECT  0.245 0.545 0.495 1.365 ;
        RECT  2.650 2.380 3.845 2.780 ;
        RECT  2.405 2.380 2.650 3.290 ;
        RECT  1.210 2.380 2.405 2.780 ;
        RECT  0.965 2.380 1.210 3.290 ;
        RECT  11.775 0.485 12.015 1.320 ;
        RECT  6.255 0.485 11.775 0.715 ;
        RECT  6.005 0.485 6.255 1.365 ;
        RECT  4.815 1.070 6.005 1.365 ;
    END
END CKND2D8BWP7T

MACRO CKND3BWP7T
    CLASS CORE ;
    FOREIGN CKND3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.9192 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 2.190 3.070 3.415 ;
        RECT  2.830 1.030 2.970 3.415 ;
        RECT  2.215 1.030 2.830 2.540 ;
        RECT  2.070 0.540 2.215 2.540 ;
        RECT  1.960 0.540 2.070 1.360 ;
        RECT  1.550 2.190 2.070 2.540 ;
        RECT  1.310 2.190 1.550 3.415 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.0233 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.480 1.655 1.700 1.895 ;
        RECT  0.140 0.960 0.480 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.050 -0.235 3.360 0.235 ;
        RECT  2.670 -0.235 3.050 0.785 ;
        RECT  1.550 -0.235 2.670 0.235 ;
        RECT  1.170 -0.235 1.550 1.210 ;
        RECT  0.000 -0.235 1.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 3.685 3.360 4.155 ;
        RECT  1.990 2.780 2.370 4.155 ;
        RECT  0.900 3.685 1.990 4.155 ;
        RECT  0.520 2.500 0.900 4.155 ;
        RECT  0.000 3.685 0.520 4.155 ;
        END
    END VDD
END CKND3BWP7T

MACRO CKND4BWP7T
    CLASS CORE ;
    FOREIGN CKND4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.2496 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 2.200 2.790 3.380 ;
        RECT  2.485 0.540 2.730 1.420 ;
        RECT  2.410 2.200 2.550 2.550 ;
        RECT  2.410 1.070 2.485 1.420 ;
        RECT  1.510 1.070 2.410 2.550 ;
        RECT  1.270 1.070 1.510 1.420 ;
        RECT  1.270 2.200 1.510 2.550 ;
        RECT  1.030 0.510 1.270 1.420 ;
        RECT  1.030 2.200 1.270 3.380 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.3644 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.705 1.200 1.950 ;
        RECT  0.140 0.905 0.470 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 -0.235 3.920 0.235 ;
        RECT  3.200 -0.235 3.580 0.835 ;
        RECT  2.060 -0.235 3.200 0.235 ;
        RECT  1.680 -0.235 2.060 0.790 ;
        RECT  0.000 -0.235 1.680 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 3.685 3.920 4.155 ;
        RECT  3.200 2.300 3.580 4.155 ;
        RECT  2.100 3.685 3.200 4.155 ;
        RECT  1.720 2.780 2.100 4.155 ;
        RECT  0.620 3.685 1.720 4.155 ;
        RECT  0.240 2.510 0.620 4.155 ;
        RECT  0.000 3.685 0.240 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.610 2.200 2.790 3.380 ;
        RECT  2.610 0.540 2.730 1.420 ;
        RECT  1.270 1.070 1.310 1.420 ;
        RECT  1.270 2.200 1.310 2.550 ;
        RECT  1.030 0.510 1.270 1.420 ;
        RECT  1.030 2.200 1.270 3.380 ;
    END
END CKND4BWP7T

MACRO CKND6BWP7T
    CLASS CORE ;
    FOREIGN CKND6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0726 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.845 0.565 4.090 1.420 ;
        RECT  3.850 2.200 4.090 3.410 ;
        RECT  2.970 2.200 3.850 2.550 ;
        RECT  2.970 1.070 3.845 1.420 ;
        RECT  2.650 1.070 2.970 2.550 ;
        RECT  2.410 0.565 2.650 3.410 ;
        RECT  2.405 0.565 2.410 2.550 ;
        RECT  2.070 1.070 2.405 2.550 ;
        RECT  1.210 2.200 2.070 2.550 ;
        RECT  0.970 2.200 1.210 3.410 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 2.0484 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.645 1.650 1.890 ;
        RECT  0.450 0.905 0.470 1.890 ;
        RECT  0.140 0.905 0.450 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 -0.235 5.040 0.235 ;
        RECT  4.500 -0.235 4.880 0.875 ;
        RECT  3.440 -0.235 4.500 0.235 ;
        RECT  3.060 -0.235 3.440 0.790 ;
        RECT  1.840 -0.235 3.060 0.235 ;
        RECT  1.590 -0.235 1.840 0.925 ;
        RECT  0.000 -0.235 1.590 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 3.685 5.040 4.155 ;
        RECT  4.500 2.300 4.880 4.155 ;
        RECT  3.440 3.685 4.500 4.155 ;
        RECT  3.060 2.780 3.440 4.155 ;
        RECT  2.000 3.685 3.060 4.155 ;
        RECT  1.620 2.780 2.000 4.155 ;
        RECT  0.560 3.685 1.620 4.155 ;
        RECT  0.180 2.560 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.845 0.565 4.090 1.420 ;
        RECT  3.850 2.200 4.090 3.410 ;
        RECT  3.170 2.200 3.850 2.550 ;
        RECT  3.170 1.070 3.845 1.420 ;
        RECT  1.210 2.200 1.870 2.550 ;
        RECT  0.970 2.200 1.210 3.410 ;
    END
END CKND6BWP7T

MACRO CKND8BWP7T
    CLASS CORE ;
    FOREIGN CKND8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 4.0932 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.285 0.515 5.530 1.420 ;
        RECT  5.290 2.150 5.530 3.405 ;
        RECT  4.090 2.150 5.290 2.550 ;
        RECT  4.090 1.020 5.285 1.420 ;
        RECT  3.850 0.515 4.090 3.405 ;
        RECT  3.845 0.515 3.850 2.550 ;
        RECT  3.190 1.020 3.845 2.550 ;
        RECT  2.650 1.020 3.190 1.420 ;
        RECT  2.650 2.150 3.190 2.550 ;
        RECT  2.405 0.515 2.650 1.420 ;
        RECT  2.410 2.150 2.650 3.405 ;
        RECT  1.210 2.150 2.410 2.550 ;
        RECT  0.970 2.150 1.210 3.405 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 2.7288 ;
        ANTENNADIFFAREA 0.2037 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.650 2.595 1.895 ;
        RECT  0.450 0.905 0.470 1.895 ;
        RECT  0.140 0.905 0.450 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.320 -0.235 6.720 0.235 ;
        RECT  5.940 -0.235 6.320 0.815 ;
        RECT  4.880 -0.235 5.940 0.235 ;
        RECT  4.500 -0.235 4.880 0.790 ;
        RECT  3.440 -0.235 4.500 0.235 ;
        RECT  3.060 -0.235 3.440 0.790 ;
        RECT  1.935 -0.235 3.060 0.235 ;
        RECT  1.685 -0.235 1.935 0.880 ;
        RECT  0.000 -0.235 1.685 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.320 3.685 6.720 4.155 ;
        RECT  5.940 2.300 6.320 4.155 ;
        RECT  4.880 3.685 5.940 4.155 ;
        RECT  4.500 2.780 4.880 4.155 ;
        RECT  3.440 3.685 4.500 4.155 ;
        RECT  3.060 2.780 3.440 4.155 ;
        RECT  2.000 3.685 3.060 4.155 ;
        RECT  1.620 2.780 2.000 4.155 ;
        RECT  0.560 3.685 1.620 4.155 ;
        RECT  0.180 2.560 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.285 0.515 5.530 1.420 ;
        RECT  5.290 2.150 5.530 3.405 ;
        RECT  4.290 2.150 5.290 2.550 ;
        RECT  4.290 1.020 5.285 1.420 ;
        RECT  2.650 1.020 2.990 1.420 ;
        RECT  2.650 2.150 2.990 2.550 ;
        RECT  2.405 0.515 2.650 1.420 ;
        RECT  2.410 2.150 2.650 3.405 ;
        RECT  1.210 2.150 2.410 2.550 ;
        RECT  0.970 2.150 1.210 3.405 ;
    END
END CKND8BWP7T

MACRO CKXOR2D0BWP7T
    CLASS CORE ;
    FOREIGN CKXOR2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.6240 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.810 0.480 4.900 2.845 ;
        RECT  4.620 0.480 4.810 3.130 ;
        RECT  4.570 0.480 4.620 0.820 ;
        RECT  4.570 2.575 4.620 3.130 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2448 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 1.210 3.830 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.5661 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 -0.235 5.040 0.235 ;
        RECT  3.780 -0.235 4.160 0.770 ;
        RECT  1.185 -0.235 3.780 0.235 ;
        RECT  0.955 -0.235 1.185 0.820 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 3.685 5.040 4.155 ;
        RECT  3.780 3.235 4.160 4.155 ;
        RECT  1.300 3.685 3.780 4.155 ;
        RECT  0.920 2.875 1.300 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.340 1.610 4.390 1.950 ;
        RECT  4.110 1.610 4.340 3.005 ;
        RECT  2.750 2.775 4.110 3.005 ;
        RECT  3.210 0.465 3.345 0.820 ;
        RECT  3.210 2.300 3.330 2.530 ;
        RECT  2.980 0.465 3.210 2.530 ;
        RECT  1.935 0.465 2.980 0.695 ;
        RECT  2.520 0.925 2.750 3.005 ;
        RECT  2.515 0.925 2.520 2.720 ;
        RECT  2.300 0.925 2.515 1.155 ;
        RECT  2.305 2.380 2.515 2.720 ;
        RECT  2.075 1.625 2.285 1.965 ;
        RECT  1.845 1.625 2.075 2.645 ;
        RECT  1.705 0.465 1.935 1.360 ;
        RECT  0.465 2.410 1.845 2.645 ;
        RECT  1.615 1.130 1.705 1.360 ;
        RECT  1.385 1.130 1.615 1.945 ;
        RECT  0.235 0.480 0.465 2.645 ;
    END
END CKXOR2D0BWP7T

MACRO CKXOR2D1BWP7T
    CLASS CORE ;
    FOREIGN CKXOR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.0416 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.810 0.480 4.900 2.805 ;
        RECT  4.620 0.480 4.810 3.455 ;
        RECT  4.570 0.480 4.620 0.820 ;
        RECT  4.570 2.535 4.620 3.455 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 1.210 3.830 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.5661 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 -0.235 5.040 0.235 ;
        RECT  3.780 -0.235 4.160 0.770 ;
        RECT  1.185 -0.235 3.780 0.235 ;
        RECT  0.955 -0.235 1.185 0.820 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 3.685 5.040 4.155 ;
        RECT  3.780 3.220 4.160 4.155 ;
        RECT  1.300 3.685 3.780 4.155 ;
        RECT  0.920 3.010 1.300 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.340 1.610 4.390 1.950 ;
        RECT  4.110 1.610 4.340 2.990 ;
        RECT  2.750 2.760 4.110 2.990 ;
        RECT  3.210 0.465 3.345 0.820 ;
        RECT  3.210 2.300 3.330 2.530 ;
        RECT  2.980 0.465 3.210 2.530 ;
        RECT  1.935 0.465 2.980 0.695 ;
        RECT  2.520 0.925 2.750 2.990 ;
        RECT  2.515 0.925 2.520 2.720 ;
        RECT  2.300 0.925 2.515 1.155 ;
        RECT  2.305 2.380 2.515 2.720 ;
        RECT  2.075 1.625 2.285 1.965 ;
        RECT  1.845 1.625 2.075 2.780 ;
        RECT  1.705 0.465 1.935 1.360 ;
        RECT  0.465 2.545 1.845 2.780 ;
        RECT  1.615 1.130 1.705 1.360 ;
        RECT  1.385 1.130 1.615 1.945 ;
        RECT  0.235 0.480 0.465 2.780 ;
    END
END CKXOR2D1BWP7T

MACRO CKXOR2D2BWP7T
    CLASS CORE ;
    FOREIGN CKXOR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 0.695 6.020 3.190 ;
        RECT  4.880 0.695 5.740 0.925 ;
        RECT  4.815 2.960 5.740 3.190 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.3240 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 1.770 4.900 2.150 ;
        RECT  3.850 1.605 4.140 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.5985 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 -0.235 6.160 0.235 ;
        RECT  5.640 -0.235 5.980 0.465 ;
        RECT  4.410 -0.235 5.640 0.235 ;
        RECT  4.175 -0.235 4.410 0.520 ;
        RECT  1.240 -0.235 4.175 0.235 ;
        RECT  0.900 -0.235 1.240 0.730 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 3.685 6.160 4.155 ;
        RECT  5.640 3.450 5.980 4.155 ;
        RECT  4.480 3.685 5.640 4.155 ;
        RECT  4.100 3.455 4.480 4.155 ;
        RECT  1.280 3.685 4.100 4.155 ;
        RECT  0.920 3.455 1.280 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.160 1.155 5.390 2.730 ;
        RECT  4.465 1.155 5.160 1.385 ;
        RECT  4.190 2.500 5.160 2.730 ;
        RECT  4.235 0.925 4.465 1.385 ;
        RECT  3.945 0.925 4.235 1.155 ;
        RECT  3.960 2.500 4.190 3.225 ;
        RECT  2.250 2.995 3.960 3.225 ;
        RECT  3.715 0.465 3.945 1.155 ;
        RECT  2.300 0.465 3.715 0.695 ;
        RECT  3.400 1.390 3.495 2.700 ;
        RECT  3.265 0.925 3.400 2.700 ;
        RECT  3.170 0.925 3.265 1.620 ;
        RECT  3.145 2.470 3.265 2.700 ;
        RECT  1.615 0.925 3.170 1.155 ;
        RECT  2.745 1.895 3.035 2.235 ;
        RECT  2.515 1.895 2.745 2.645 ;
        RECT  2.010 2.415 2.515 2.645 ;
        RECT  2.075 1.545 2.285 1.885 ;
        RECT  1.845 1.545 2.075 2.160 ;
        RECT  1.780 2.415 2.010 3.115 ;
        RECT  1.445 1.925 1.845 2.160 ;
        RECT  0.705 2.885 1.780 3.115 ;
        RECT  1.385 0.925 1.615 1.695 ;
        RECT  1.210 1.925 1.445 2.655 ;
        RECT  0.465 2.420 1.210 2.655 ;
        RECT  0.475 2.885 0.705 3.305 ;
        RECT  0.235 0.480 0.465 2.655 ;
    END
END CKXOR2D2BWP7T

MACRO CKXOR2D4BWP7T
    CLASS CORE ;
    FOREIGN CKXOR2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.1276 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.135 0.580 11.370 3.220 ;
        RECT  10.470 1.140 11.135 2.505 ;
        RECT  9.930 1.140 10.470 1.430 ;
        RECT  9.930 2.155 10.470 2.505 ;
        RECT  9.690 0.655 9.930 1.430 ;
        RECT  9.695 2.155 9.930 3.220 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 1.0098 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.730 7.755 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8883 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.515 2.295 1.855 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.160 -0.235 12.320 0.235 ;
        RECT  11.780 -0.235 12.160 0.955 ;
        RECT  10.720 -0.235 11.780 0.235 ;
        RECT  10.340 -0.235 10.720 0.885 ;
        RECT  9.205 -0.235 10.340 0.235 ;
        RECT  8.975 -0.235 9.205 0.935 ;
        RECT  7.295 -0.235 8.975 0.235 ;
        RECT  7.065 -0.235 7.295 0.935 ;
        RECT  1.945 -0.235 7.065 0.235 ;
        RECT  1.715 -0.235 1.945 0.520 ;
        RECT  0.465 -0.235 1.715 0.235 ;
        RECT  0.235 -0.235 0.465 0.980 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.160 3.685 12.320 4.155 ;
        RECT  11.780 2.305 12.160 4.155 ;
        RECT  10.720 3.685 11.780 4.155 ;
        RECT  10.340 2.780 10.720 4.155 ;
        RECT  9.275 3.685 10.340 4.155 ;
        RECT  8.895 2.300 9.275 4.155 ;
        RECT  7.840 3.685 8.895 4.155 ;
        RECT  7.460 3.055 7.840 4.155 ;
        RECT  1.905 3.685 7.460 4.155 ;
        RECT  1.620 3.040 1.905 4.155 ;
        RECT  0.540 3.685 1.620 4.155 ;
        RECT  0.160 2.310 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.930 1.140 10.270 1.430 ;
        RECT  9.930 2.155 10.270 2.505 ;
        RECT  9.690 0.655 9.930 1.430 ;
        RECT  9.695 2.155 9.930 3.220 ;
        RECT  8.745 1.660 10.210 1.895 ;
        RECT  8.515 0.465 8.745 1.895 ;
        RECT  7.755 0.465 8.515 0.695 ;
        RECT  8.250 2.440 8.490 3.360 ;
        RECT  8.235 2.440 8.250 2.690 ;
        RECT  8.005 0.925 8.235 2.690 ;
        RECT  7.050 2.440 8.005 2.690 ;
        RECT  7.525 0.465 7.755 1.490 ;
        RECT  6.520 1.250 7.525 1.490 ;
        RECT  6.810 2.440 7.050 3.455 ;
        RECT  5.635 3.215 6.810 3.455 ;
        RECT  6.500 0.465 6.520 1.490 ;
        RECT  6.350 0.465 6.500 2.780 ;
        RECT  6.260 0.465 6.350 2.935 ;
        RECT  5.065 0.465 6.260 0.695 ;
        RECT  6.110 2.490 6.260 2.935 ;
        RECT  5.635 0.925 5.840 1.155 ;
        RECT  5.390 0.925 5.635 3.455 ;
        RECT  2.365 3.225 5.390 3.455 ;
        RECT  4.830 0.465 5.065 2.995 ;
        RECT  4.670 2.520 4.830 2.995 ;
        RECT  3.565 2.765 4.670 2.995 ;
        RECT  4.110 0.465 4.350 2.440 ;
        RECT  2.405 0.465 4.110 0.695 ;
        RECT  3.900 2.205 4.110 2.440 ;
        RECT  3.565 0.925 3.675 1.155 ;
        RECT  3.325 0.925 3.565 2.995 ;
        RECT  3.075 2.760 3.325 2.995 ;
        RECT  2.975 1.595 3.095 1.935 ;
        RECT  2.790 0.925 2.975 1.935 ;
        RECT  2.635 0.925 2.790 2.490 ;
        RECT  2.555 1.540 2.635 2.490 ;
        RECT  2.175 0.465 2.405 0.980 ;
        RECT  2.325 2.705 2.365 3.455 ;
        RECT  2.135 2.480 2.325 3.455 ;
        RECT  1.240 0.750 2.175 0.980 ;
        RECT  2.095 2.480 2.135 2.885 ;
        RECT  1.570 2.480 2.095 2.710 ;
        RECT  1.290 1.335 1.570 2.710 ;
        RECT  1.040 0.720 1.240 0.980 ;
        RECT  1.040 2.960 1.240 3.200 ;
        RECT  0.810 0.720 1.040 3.200 ;
    END
END CKXOR2D4BWP7T

MACRO DCAP16BWP7T
    CLASS CORE ;
    FOREIGN DCAP16BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.080 -0.235 8.960 0.235 ;
        RECT  7.700 -0.235 8.080 0.785 ;
        RECT  6.565 -0.235 7.700 0.235 ;
        RECT  6.185 -0.235 6.565 1.215 ;
        RECT  5.060 -0.235 6.185 0.235 ;
        RECT  4.680 -0.235 5.060 1.215 ;
        RECT  3.555 -0.235 4.680 0.235 ;
        RECT  3.175 -0.235 3.555 1.215 ;
        RECT  2.050 -0.235 3.175 0.235 ;
        RECT  1.670 -0.235 2.050 1.215 ;
        RECT  0.545 -0.235 1.670 0.235 ;
        RECT  0.165 -0.235 0.545 1.215 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.085 3.685 8.960 4.155 ;
        RECT  7.705 2.655 8.085 4.155 ;
        RECT  6.565 3.685 7.705 4.155 ;
        RECT  6.185 2.680 6.565 4.155 ;
        RECT  5.060 3.685 6.185 4.155 ;
        RECT  4.680 2.680 5.060 4.155 ;
        RECT  3.555 3.685 4.680 4.155 ;
        RECT  3.175 2.680 3.555 4.155 ;
        RECT  2.050 3.685 3.175 4.155 ;
        RECT  1.670 2.595 2.050 4.155 ;
        RECT  0.560 3.685 1.670 4.155 ;
        RECT  0.180 2.595 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.495 1.485 8.740 3.410 ;
        RECT  8.495 0.660 8.725 1.255 ;
        RECT  7.765 1.015 8.495 1.255 ;
        RECT  7.535 1.015 7.765 2.225 ;
        RECT  6.765 1.995 7.535 2.225 ;
    END
END DCAP16BWP7T

MACRO DCAP32BWP7T
    CLASS CORE ;
    FOREIGN DCAP32BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.035 -0.235 17.920 0.235 ;
        RECT  16.655 -0.235 17.035 0.780 ;
        RECT  15.430 -0.235 16.655 0.235 ;
        RECT  15.050 -0.235 15.430 1.230 ;
        RECT  13.855 -0.235 15.050 0.235 ;
        RECT  13.475 -0.235 13.855 1.230 ;
        RECT  12.280 -0.235 13.475 0.235 ;
        RECT  11.900 -0.235 12.280 1.230 ;
        RECT  10.705 -0.235 11.900 0.235 ;
        RECT  10.325 -0.235 10.705 1.230 ;
        RECT  9.135 -0.235 10.325 0.235 ;
        RECT  8.755 -0.235 9.135 1.220 ;
        RECT  7.560 -0.235 8.755 0.235 ;
        RECT  7.180 -0.235 7.560 1.220 ;
        RECT  5.985 -0.235 7.180 0.235 ;
        RECT  5.605 -0.235 5.985 1.220 ;
        RECT  4.410 -0.235 5.605 0.235 ;
        RECT  4.030 -0.235 4.410 1.220 ;
        RECT  2.835 -0.235 4.030 0.235 ;
        RECT  2.455 -0.235 2.835 1.220 ;
        RECT  1.240 -0.235 2.455 0.235 ;
        RECT  0.860 -0.235 1.240 0.780 ;
        RECT  0.000 -0.235 0.860 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.000 3.685 17.920 4.155 ;
        RECT  16.620 2.650 17.000 4.155 ;
        RECT  15.425 3.685 16.620 4.155 ;
        RECT  15.045 2.650 15.425 4.155 ;
        RECT  13.850 3.685 15.045 4.155 ;
        RECT  13.470 2.460 13.850 4.155 ;
        RECT  12.275 3.685 13.470 4.155 ;
        RECT  11.895 2.460 12.275 4.155 ;
        RECT  10.700 3.685 11.895 4.155 ;
        RECT  10.320 2.460 10.700 4.155 ;
        RECT  9.125 3.685 10.320 4.155 ;
        RECT  8.745 2.460 9.125 4.155 ;
        RECT  7.550 3.685 8.745 4.155 ;
        RECT  7.170 2.440 7.550 4.155 ;
        RECT  5.975 3.685 7.170 4.155 ;
        RECT  5.595 2.440 5.975 4.155 ;
        RECT  4.400 3.685 5.595 4.155 ;
        RECT  4.020 2.440 4.400 4.155 ;
        RECT  2.825 3.685 4.020 4.155 ;
        RECT  2.445 2.630 2.825 4.155 ;
        RECT  1.250 3.685 2.445 4.155 ;
        RECT  0.870 2.630 1.250 4.155 ;
        RECT  0.000 3.685 0.870 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.455 1.485 17.700 3.405 ;
        RECT  17.455 0.680 17.685 1.255 ;
        RECT  17.085 1.015 17.455 1.255 ;
        RECT  16.845 1.015 17.085 2.225 ;
        RECT  16.275 1.995 16.845 2.225 ;
        RECT  1.280 1.995 1.910 2.225 ;
        RECT  1.040 1.015 1.280 2.225 ;
        RECT  0.465 1.015 1.040 1.255 ;
        RECT  0.235 0.635 0.465 1.255 ;
        RECT  0.220 1.485 0.465 3.385 ;
    END
END DCAP32BWP7T

MACRO DCAP4BWP7T
    CLASS CORE ;
    FOREIGN DCAP4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.360 -0.235 2.240 0.235 ;
        RECT  0.980 -0.235 1.360 1.200 ;
        RECT  0.545 -0.235 0.980 0.235 ;
        RECT  0.165 -0.235 0.545 1.200 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.375 3.685 2.240 4.155 ;
        RECT  0.995 3.050 1.375 4.155 ;
        RECT  0.550 3.685 0.995 4.155 ;
        RECT  0.170 2.635 0.550 4.155 ;
        RECT  0.000 3.685 0.170 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.775 0.495 2.020 2.265 ;
        RECT  1.775 2.580 2.005 3.390 ;
        RECT  1.040 2.580 1.775 2.820 ;
        RECT  0.800 1.540 1.040 2.820 ;
        RECT  0.165 1.540 0.800 1.770 ;
    END
END DCAP4BWP7T

MACRO DCAP64BWP7T
    CLASS CORE ;
    FOREIGN DCAP64BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.840 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  34.955 -0.235 35.840 0.235 ;
        RECT  34.575 -0.235 34.955 0.760 ;
        RECT  33.390 -0.235 34.575 0.235 ;
        RECT  33.010 -0.235 33.390 1.220 ;
        RECT  31.860 -0.235 33.010 0.235 ;
        RECT  31.480 -0.235 31.860 1.220 ;
        RECT  30.330 -0.235 31.480 0.235 ;
        RECT  29.950 -0.235 30.330 1.220 ;
        RECT  28.800 -0.235 29.950 0.235 ;
        RECT  28.420 -0.235 28.800 1.220 ;
        RECT  27.270 -0.235 28.420 0.235 ;
        RECT  26.890 -0.235 27.270 1.220 ;
        RECT  25.740 -0.235 26.890 0.235 ;
        RECT  25.360 -0.235 25.740 1.220 ;
        RECT  24.210 -0.235 25.360 0.235 ;
        RECT  23.830 -0.235 24.210 1.220 ;
        RECT  22.680 -0.235 23.830 0.235 ;
        RECT  22.300 -0.235 22.680 1.220 ;
        RECT  21.150 -0.235 22.300 0.235 ;
        RECT  20.770 -0.235 21.150 1.220 ;
        RECT  19.620 -0.235 20.770 0.235 ;
        RECT  19.240 -0.235 19.620 1.220 ;
        RECT  18.090 -0.235 19.240 0.235 ;
        RECT  17.710 -0.235 18.090 1.220 ;
        RECT  16.560 -0.235 17.710 0.235 ;
        RECT  16.180 -0.235 16.560 1.220 ;
        RECT  15.030 -0.235 16.180 0.235 ;
        RECT  14.650 -0.235 15.030 1.220 ;
        RECT  13.500 -0.235 14.650 0.235 ;
        RECT  13.120 -0.235 13.500 1.220 ;
        RECT  11.970 -0.235 13.120 0.235 ;
        RECT  11.590 -0.235 11.970 1.220 ;
        RECT  10.440 -0.235 11.590 0.235 ;
        RECT  10.060 -0.235 10.440 1.220 ;
        RECT  8.910 -0.235 10.060 0.235 ;
        RECT  8.530 -0.235 8.910 1.220 ;
        RECT  7.380 -0.235 8.530 0.235 ;
        RECT  7.000 -0.235 7.380 1.220 ;
        RECT  5.850 -0.235 7.000 0.235 ;
        RECT  5.470 -0.235 5.850 1.220 ;
        RECT  4.320 -0.235 5.470 0.235 ;
        RECT  3.940 -0.235 4.320 1.220 ;
        RECT  2.790 -0.235 3.940 0.235 ;
        RECT  2.410 -0.235 2.790 1.220 ;
        RECT  1.240 -0.235 2.410 0.235 ;
        RECT  0.860 -0.235 1.240 0.780 ;
        RECT  0.000 -0.235 0.860 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  34.950 3.685 35.840 4.155 ;
        RECT  34.570 2.650 34.950 4.155 ;
        RECT  33.380 3.685 34.570 4.155 ;
        RECT  33.000 2.650 33.380 4.155 ;
        RECT  31.850 3.685 33.000 4.155 ;
        RECT  31.470 2.650 31.850 4.155 ;
        RECT  30.320 3.685 31.470 4.155 ;
        RECT  29.940 2.650 30.320 4.155 ;
        RECT  28.790 3.685 29.940 4.155 ;
        RECT  28.410 2.650 28.790 4.155 ;
        RECT  27.260 3.685 28.410 4.155 ;
        RECT  26.880 2.650 27.260 4.155 ;
        RECT  25.730 3.685 26.880 4.155 ;
        RECT  25.350 2.650 25.730 4.155 ;
        RECT  24.200 3.685 25.350 4.155 ;
        RECT  23.820 2.650 24.200 4.155 ;
        RECT  22.670 3.685 23.820 4.155 ;
        RECT  22.290 2.650 22.670 4.155 ;
        RECT  21.140 3.685 22.290 4.155 ;
        RECT  20.760 2.650 21.140 4.155 ;
        RECT  19.610 3.685 20.760 4.155 ;
        RECT  19.230 2.650 19.610 4.155 ;
        RECT  18.080 3.685 19.230 4.155 ;
        RECT  17.700 2.650 18.080 4.155 ;
        RECT  16.550 3.685 17.700 4.155 ;
        RECT  16.170 2.650 16.550 4.155 ;
        RECT  15.020 3.685 16.170 4.155 ;
        RECT  14.640 2.650 15.020 4.155 ;
        RECT  13.490 3.685 14.640 4.155 ;
        RECT  13.110 2.650 13.490 4.155 ;
        RECT  11.960 3.685 13.110 4.155 ;
        RECT  11.580 2.650 11.960 4.155 ;
        RECT  10.430 3.685 11.580 4.155 ;
        RECT  10.050 2.650 10.430 4.155 ;
        RECT  8.900 3.685 10.050 4.155 ;
        RECT  8.520 2.650 8.900 4.155 ;
        RECT  7.370 3.685 8.520 4.155 ;
        RECT  6.990 2.630 7.370 4.155 ;
        RECT  5.840 3.685 6.990 4.155 ;
        RECT  5.460 2.630 5.840 4.155 ;
        RECT  4.310 3.685 5.460 4.155 ;
        RECT  3.930 2.630 4.310 4.155 ;
        RECT  2.780 3.685 3.930 4.155 ;
        RECT  2.400 2.630 2.780 4.155 ;
        RECT  1.250 3.685 2.400 4.155 ;
        RECT  0.870 2.630 1.250 4.155 ;
        RECT  0.000 3.685 0.870 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  35.375 1.485 35.620 3.405 ;
        RECT  35.375 0.690 35.605 1.230 ;
        RECT  34.915 0.990 35.375 1.230 ;
        RECT  34.675 0.990 34.915 2.225 ;
        RECT  34.105 1.995 34.675 2.225 ;
        RECT  1.280 1.995 1.910 2.225 ;
        RECT  1.040 1.015 1.280 2.225 ;
        RECT  0.465 1.015 1.040 1.255 ;
        RECT  0.235 0.695 0.465 1.255 ;
        RECT  0.220 1.485 0.465 3.385 ;
    END
END DCAP64BWP7T

MACRO DCAP8BWP7T
    CLASS CORE ;
    FOREIGN DCAP8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.600 -0.235 4.480 0.235 ;
        RECT  3.220 -0.235 3.600 0.700 ;
        RECT  2.070 -0.235 3.220 0.235 ;
        RECT  1.690 -0.235 2.070 1.165 ;
        RECT  0.540 -0.235 1.690 0.235 ;
        RECT  0.160 -0.235 0.540 1.165 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.600 3.685 4.480 4.155 ;
        RECT  3.220 2.510 3.600 4.155 ;
        RECT  2.050 3.685 3.220 4.155 ;
        RECT  1.710 2.510 2.050 4.155 ;
        RECT  0.520 3.685 1.710 4.155 ;
        RECT  0.180 2.510 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.015 0.620 4.245 1.170 ;
        RECT  4.015 1.430 4.245 3.265 ;
        RECT  3.625 0.930 4.015 1.170 ;
        RECT  3.385 0.930 3.625 2.145 ;
        RECT  2.645 1.915 3.385 2.145 ;
    END
END DCAP8BWP7T

MACRO DCAPBWP7T
    CLASS CORE ;
    FOREIGN DCAPBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.640 -0.235 1.680 0.235 ;
        RECT  0.300 -0.235 0.640 0.765 ;
        RECT  0.000 -0.235 0.300 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.560 3.685 1.680 4.155 ;
        RECT  0.220 2.645 0.560 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.290 1.560 1.490 1.790 ;
        RECT  1.140 0.470 1.370 1.280 ;
        RECT  1.060 1.560 1.290 3.450 ;
        RECT  0.455 1.050 1.140 1.280 ;
        RECT  0.225 1.050 0.455 2.065 ;
    END
END DCAPBWP7T

MACRO DEL015BWP7T
    CLASS CORE ;
    FOREIGN DEL015BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.7584 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.510 2.100 3.360 ;
        RECT  1.625 0.510 1.820 0.740 ;
        RECT  1.625 3.130 1.820 3.360 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.130 1.770 0.980 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 -0.235 2.240 0.235 ;
        RECT  0.875 -0.235 1.290 0.720 ;
        RECT  0.000 -0.235 0.875 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 3.685 2.240 4.155 ;
        RECT  0.890 3.040 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.355 1.310 1.585 2.765 ;
        RECT  0.470 1.310 1.355 1.540 ;
        RECT  0.470 2.525 1.355 2.765 ;
        RECT  0.240 0.495 0.470 1.540 ;
        RECT  0.240 2.525 0.470 3.390 ;
    END
END DEL015BWP7T

MACRO DEL01BWP7T
    CLASS CORE ;
    FOREIGN DEL01BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.585 2.100 3.360 ;
        RECT  1.625 0.585 1.820 0.815 ;
        RECT  1.625 3.130 1.820 3.360 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.130 1.770 0.980 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 -0.235 2.240 0.235 ;
        RECT  0.875 -0.235 1.290 0.780 ;
        RECT  0.000 -0.235 0.875 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 3.685 2.240 4.155 ;
        RECT  0.890 3.040 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.355 1.135 1.585 2.735 ;
        RECT  0.470 1.135 1.355 1.365 ;
        RECT  0.470 2.495 1.355 2.735 ;
        RECT  0.240 0.590 0.470 1.365 ;
        RECT  0.240 2.495 0.470 3.390 ;
    END
END DEL01BWP7T

MACRO DEL02BWP7T
    CLASS CORE ;
    FOREIGN DEL02BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5184 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.780 2.100 3.360 ;
        RECT  1.625 0.780 1.820 1.010 ;
        RECT  1.625 3.130 1.820 3.360 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2124 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.130 1.770 0.980 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 -0.235 2.240 0.235 ;
        RECT  0.875 -0.235 1.290 1.010 ;
        RECT  0.000 -0.235 0.875 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.295 3.685 2.240 4.155 ;
        RECT  0.890 3.010 1.295 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.355 1.310 1.585 2.765 ;
        RECT  0.470 1.310 1.355 1.540 ;
        RECT  0.470 2.525 1.355 2.765 ;
        RECT  0.240 0.565 0.470 1.540 ;
        RECT  0.240 2.525 0.470 3.335 ;
    END
END DEL02BWP7T

MACRO DEL0BWP7T
    CLASS CORE ;
    FOREIGN DEL0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.465 4.340 3.335 ;
        RECT  3.960 0.465 4.060 0.695 ;
        RECT  3.960 2.635 4.060 3.335 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.595 -0.235 4.480 0.235 ;
        RECT  3.185 -0.235 3.595 0.775 ;
        RECT  1.285 -0.235 3.185 0.235 ;
        RECT  0.875 -0.235 1.285 0.670 ;
        RECT  0.000 -0.235 0.875 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 3.685 4.480 4.155 ;
        RECT  3.225 3.110 3.590 4.155 ;
        RECT  1.270 3.685 3.225 4.155 ;
        RECT  0.890 3.105 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.485 1.190 3.715 2.725 ;
        RECT  2.705 1.190 3.485 1.430 ;
        RECT  2.705 2.495 3.485 2.725 ;
        RECT  2.210 1.765 3.085 1.995 ;
        RECT  2.475 0.490 2.705 1.430 ;
        RECT  2.475 2.495 2.705 3.330 ;
        RECT  1.980 0.545 2.210 3.170 ;
        RECT  1.720 0.545 1.980 0.775 ;
        RECT  1.685 2.930 1.980 3.170 ;
        RECT  1.435 1.250 1.665 2.030 ;
        RECT  0.465 1.250 1.435 1.530 ;
        RECT  0.235 0.465 0.465 3.265 ;
    END
END DEL0BWP7T

MACRO DEL1BWP7T
    CLASS CORE ;
    FOREIGN DEL1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.325 0.655 5.460 2.810 ;
        RECT  5.180 0.655 5.325 3.390 ;
        RECT  5.040 0.655 5.180 0.885 ;
        RECT  5.095 2.580 5.180 3.390 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.750 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.685 -0.235 5.600 0.235 ;
        RECT  4.305 -0.235 4.685 0.935 ;
        RECT  1.270 -0.235 4.305 0.235 ;
        RECT  0.890 -0.235 1.270 0.890 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.685 3.685 5.600 4.155 ;
        RECT  4.305 2.770 4.685 4.155 ;
        RECT  1.270 3.685 4.305 4.155 ;
        RECT  0.890 3.025 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.615 1.165 4.845 2.395 ;
        RECT  3.245 1.165 4.615 1.405 ;
        RECT  3.245 2.115 4.615 2.395 ;
        RECT  2.545 1.655 3.915 1.885 ;
        RECT  3.015 0.650 3.245 1.405 ;
        RECT  3.015 2.115 3.245 3.290 ;
        RECT  2.315 0.790 2.545 3.370 ;
        RECT  1.585 1.175 1.815 1.945 ;
        RECT  0.465 1.175 1.585 1.455 ;
        RECT  0.235 0.595 0.465 3.310 ;
    END
END DEL1BWP7T

MACRO DEL2BWP7T
    CLASS CORE ;
    FOREIGN DEL2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.305 0.655 6.580 2.810 ;
        RECT  6.300 0.655 6.305 3.390 ;
        RECT  6.020 0.655 6.300 0.885 ;
        RECT  6.075 2.580 6.300 3.390 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 1.770 1.540 2.150 ;
        RECT  0.700 1.510 0.950 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.665 -0.235 6.720 0.235 ;
        RECT  5.285 -0.235 5.665 0.935 ;
        RECT  1.305 -0.235 5.285 0.235 ;
        RECT  0.855 -0.235 1.305 0.750 ;
        RECT  0.000 -0.235 0.855 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.665 3.685 6.720 4.155 ;
        RECT  5.285 3.160 5.665 4.155 ;
        RECT  1.270 3.685 5.285 4.155 ;
        RECT  0.890 3.110 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.595 1.165 5.825 2.395 ;
        RECT  3.795 1.165 5.595 1.405 ;
        RECT  3.795 2.150 5.595 2.395 ;
        RECT  2.975 1.655 4.905 1.885 ;
        RECT  3.565 0.650 3.795 1.405 ;
        RECT  3.565 2.150 3.795 3.425 ;
        RECT  2.745 0.465 2.975 3.280 ;
        RECT  2.005 1.030 2.235 2.145 ;
        RECT  0.465 1.030 2.005 1.280 ;
        RECT  0.235 0.465 0.465 3.390 ;
    END
END DEL2BWP7T

MACRO DEL3BWP7T
    CLASS CORE ;
    FOREIGN DEL3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.265 0.655 9.380 2.810 ;
        RECT  9.100 0.655 9.265 3.390 ;
        RECT  8.980 0.655 9.100 0.885 ;
        RECT  9.035 2.580 9.100 3.390 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.510 0.980 2.750 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.625 -0.235 9.520 0.235 ;
        RECT  8.245 -0.235 8.625 0.935 ;
        RECT  4.945 -0.235 8.245 0.235 ;
        RECT  4.565 -0.235 4.945 0.935 ;
        RECT  1.310 -0.235 4.565 0.235 ;
        RECT  0.860 -0.235 1.310 0.750 ;
        RECT  0.000 -0.235 0.860 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.625 3.685 9.520 4.155 ;
        RECT  8.245 3.000 8.625 4.155 ;
        RECT  4.960 3.685 8.245 4.155 ;
        RECT  4.555 3.250 4.960 4.155 ;
        RECT  1.270 3.685 4.555 4.155 ;
        RECT  0.890 3.110 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.555 1.165 8.785 2.395 ;
        RECT  7.055 1.165 8.555 1.405 ;
        RECT  7.055 2.115 8.555 2.395 ;
        RECT  6.355 1.655 8.070 1.885 ;
        RECT  6.825 0.650 7.055 1.405 ;
        RECT  6.825 2.115 7.055 3.295 ;
        RECT  6.125 0.650 6.355 3.400 ;
        RECT  5.365 1.775 5.860 2.115 ;
        RECT  5.115 1.165 5.365 3.020 ;
        RECT  3.375 1.165 5.115 1.405 ;
        RECT  3.375 2.775 5.115 3.020 ;
        RECT  3.730 1.655 4.070 2.355 ;
        RECT  2.675 1.655 3.730 1.935 ;
        RECT  3.145 0.650 3.375 1.405 ;
        RECT  3.145 2.775 3.375 3.350 ;
        RECT  2.445 0.465 2.675 3.315 ;
        RECT  1.665 1.025 1.895 1.880 ;
        RECT  0.465 1.025 1.665 1.255 ;
        RECT  0.235 0.465 0.465 3.390 ;
    END
END DEL3BWP7T

MACRO DEL4BWP7T
    CLASS CORE ;
    FOREIGN DEL4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.220 0.675 10.500 3.380 ;
        RECT  10.120 0.675 10.220 0.905 ;
        RECT  10.175 2.410 10.220 3.380 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.700 0.980 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.770 -0.235 10.640 0.235 ;
        RECT  9.390 -0.235 9.770 0.865 ;
        RECT  5.530 -0.235 9.390 0.235 ;
        RECT  5.150 -0.235 5.530 0.820 ;
        RECT  1.270 -0.235 5.150 0.235 ;
        RECT  0.890 -0.235 1.270 0.865 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.750 3.685 10.640 4.155 ;
        RECT  9.395 3.030 9.750 4.155 ;
        RECT  5.530 3.685 9.395 4.155 ;
        RECT  5.150 3.185 5.530 4.155 ;
        RECT  1.280 3.685 5.150 4.155 ;
        RECT  0.900 3.025 1.280 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.695 1.130 9.925 2.560 ;
        RECT  7.945 1.130 9.695 1.370 ;
        RECT  7.945 2.280 9.695 2.560 ;
        RECT  7.185 1.645 9.140 1.875 ;
        RECT  7.715 0.580 7.945 1.370 ;
        RECT  7.715 2.280 7.945 3.295 ;
        RECT  6.955 0.650 7.185 3.400 ;
        RECT  5.470 1.645 6.600 1.875 ;
        RECT  5.230 1.130 5.470 2.560 ;
        RECT  3.705 1.130 5.230 1.370 ;
        RECT  3.705 2.280 5.230 2.560 ;
        RECT  2.925 1.655 4.850 1.885 ;
        RECT  3.475 0.685 3.705 1.370 ;
        RECT  3.475 2.280 3.705 3.350 ;
        RECT  2.695 0.630 2.925 3.350 ;
        RECT  1.580 1.665 2.310 1.895 ;
        RECT  1.340 1.110 1.580 1.895 ;
        RECT  0.465 1.110 1.340 1.390 ;
        RECT  0.235 0.600 0.465 3.380 ;
    END
END DEL4BWP7T

MACRO DFCND0BWP7T
    CLASS CORE ;
    FOREIGN DFCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.340 1.200 11.620 2.560 ;
        RECT  11.205 1.200 11.340 1.430 ;
        RECT  10.970 2.330 11.340 2.560 ;
        RECT  10.975 0.605 11.205 1.430 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.410 0.605 12.740 2.715 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4158 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.725 3.385 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.700 1.540 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.455 3.225 8.345 3.455 ;
        RECT  7.225 2.730 7.455 3.455 ;
        RECT  6.290 2.730 7.225 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.980 -0.235 12.880 0.235 ;
        RECT  11.640 -0.235 11.980 0.905 ;
        RECT  8.685 -0.235 11.640 0.235 ;
        RECT  8.345 -0.235 8.685 0.465 ;
        RECT  5.570 -0.235 8.345 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  2.560 -0.235 5.230 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.915 3.685 12.880 4.155 ;
        RECT  11.575 3.455 11.915 4.155 ;
        RECT  10.810 3.685 11.575 4.155 ;
        RECT  10.470 3.455 10.810 4.155 ;
        RECT  9.280 3.685 10.470 4.155 ;
        RECT  8.940 3.190 9.280 4.155 ;
        RECT  6.995 3.685 8.940 4.155 ;
        RECT  6.655 3.190 6.995 4.155 ;
        RECT  2.385 3.685 6.655 4.155 ;
        RECT  2.045 3.455 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.935 1.600 12.165 3.020 ;
        RECT  10.720 2.790 11.935 3.020 ;
        RECT  9.165 0.465 10.740 0.695 ;
        RECT  10.490 0.990 10.720 3.020 ;
        RECT  9.695 0.990 10.490 1.220 ;
        RECT  9.995 2.510 10.490 2.740 ;
        RECT  10.005 1.565 10.235 2.280 ;
        RECT  9.345 2.050 10.005 2.280 ;
        RECT  9.765 2.510 9.995 3.375 ;
        RECT  9.465 0.990 9.695 1.820 ;
        RECT  8.680 1.590 9.465 1.820 ;
        RECT  9.115 2.050 9.345 2.960 ;
        RECT  8.935 0.465 9.165 1.220 ;
        RECT  7.915 2.730 9.115 2.960 ;
        RECT  8.405 0.990 8.935 1.220 ;
        RECT  8.405 2.270 8.690 2.500 ;
        RECT  8.175 0.990 8.405 2.500 ;
        RECT  7.435 0.990 8.175 1.220 ;
        RECT  7.685 1.615 7.915 2.960 ;
        RECT  7.140 1.615 7.685 1.845 ;
        RECT  6.910 0.985 7.140 1.845 ;
        RECT  6.505 2.270 7.060 2.500 ;
        RECT  6.715 0.985 6.910 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.075 2.460 5.735 2.690 ;
        RECT  3.845 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  3.140 0.465 4.145 0.695 ;
        RECT  1.650 2.980 3.935 3.210 ;
        RECT  3.615 0.990 3.845 2.690 ;
        RECT  3.490 0.990 3.615 1.220 ;
        RECT  3.320 2.460 3.615 2.690 ;
        RECT  2.910 0.465 3.140 1.205 ;
        RECT  2.095 0.975 2.910 1.205 ;
        RECT  1.865 0.975 2.095 2.680 ;
        RECT  1.520 0.975 1.865 1.205 ;
        RECT  1.520 2.450 1.865 2.680 ;
        RECT  1.310 2.980 1.650 3.455 ;
        RECT  0.465 2.980 1.310 3.210 ;
        RECT  0.345 0.975 0.530 1.205 ;
        RECT  0.345 2.470 0.465 3.210 ;
        RECT  0.235 0.975 0.345 3.210 ;
        RECT  0.115 0.975 0.235 2.810 ;
    END
END DFCND0BWP7T

MACRO DFCND1BWP7T
    CLASS CORE ;
    FOREIGN DFCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.8520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.340 1.075 11.620 2.560 ;
        RECT  11.205 1.075 11.340 1.305 ;
        RECT  10.970 2.330 11.340 2.560 ;
        RECT  10.975 0.480 11.205 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.410 0.470 12.740 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4158 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.725 3.385 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.700 1.540 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.455 3.225 8.345 3.455 ;
        RECT  7.225 2.730 7.455 3.455 ;
        RECT  6.290 2.730 7.225 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.980 -0.235 12.880 0.235 ;
        RECT  11.640 -0.235 11.980 0.810 ;
        RECT  8.685 -0.235 11.640 0.235 ;
        RECT  8.345 -0.235 8.685 0.465 ;
        RECT  5.570 -0.235 8.345 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  2.560 -0.235 5.230 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.915 3.685 12.880 4.155 ;
        RECT  11.575 3.455 11.915 4.155 ;
        RECT  10.810 3.685 11.575 4.155 ;
        RECT  10.470 3.455 10.810 4.155 ;
        RECT  9.280 3.685 10.470 4.155 ;
        RECT  8.940 3.190 9.280 4.155 ;
        RECT  6.995 3.685 8.940 4.155 ;
        RECT  6.655 3.190 6.995 4.155 ;
        RECT  2.385 3.685 6.655 4.155 ;
        RECT  2.045 3.455 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.935 1.600 12.165 3.020 ;
        RECT  10.720 2.790 11.935 3.020 ;
        RECT  9.165 0.465 10.740 0.695 ;
        RECT  10.490 0.990 10.720 3.020 ;
        RECT  9.695 0.990 10.490 1.220 ;
        RECT  9.995 2.565 10.490 2.795 ;
        RECT  10.005 1.565 10.235 2.260 ;
        RECT  9.345 2.030 10.005 2.260 ;
        RECT  9.765 2.565 9.995 3.375 ;
        RECT  9.465 0.990 9.695 1.760 ;
        RECT  8.680 1.530 9.465 1.760 ;
        RECT  9.115 2.030 9.345 2.960 ;
        RECT  8.935 0.465 9.165 1.220 ;
        RECT  7.915 2.730 9.115 2.960 ;
        RECT  8.405 0.990 8.935 1.220 ;
        RECT  8.405 2.270 8.690 2.500 ;
        RECT  8.175 0.990 8.405 2.500 ;
        RECT  7.435 0.990 8.175 1.220 ;
        RECT  7.685 1.615 7.915 2.960 ;
        RECT  7.140 1.615 7.685 1.845 ;
        RECT  6.910 0.985 7.140 1.845 ;
        RECT  6.505 2.270 7.060 2.500 ;
        RECT  6.715 0.985 6.910 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.075 2.460 5.735 2.690 ;
        RECT  3.845 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  3.140 0.465 4.145 0.695 ;
        RECT  1.650 2.980 3.935 3.210 ;
        RECT  3.615 0.990 3.845 2.690 ;
        RECT  3.490 0.990 3.615 1.220 ;
        RECT  3.320 2.460 3.615 2.690 ;
        RECT  2.910 0.465 3.140 1.205 ;
        RECT  2.095 0.975 2.910 1.205 ;
        RECT  1.865 0.975 2.095 2.680 ;
        RECT  1.520 0.975 1.865 1.205 ;
        RECT  1.520 2.450 1.865 2.680 ;
        RECT  1.310 2.980 1.650 3.455 ;
        RECT  0.465 2.980 1.310 3.210 ;
        RECT  0.345 0.975 0.530 1.205 ;
        RECT  0.345 2.470 0.465 3.210 ;
        RECT  0.235 0.975 0.345 3.210 ;
        RECT  0.115 0.975 0.235 2.810 ;
    END
END DFCND1BWP7T

MACRO DFCND2BWP7T
    CLASS CORE ;
    FOREIGN DFCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.880 0.465 12.225 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.605 1.055 13.860 2.690 ;
        RECT  13.580 0.465 13.605 3.310 ;
        RECT  13.370 0.465 13.580 1.285 ;
        RECT  13.375 2.460 13.580 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4158 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.725 3.385 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.700 1.540 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.455 3.225 8.355 3.455 ;
        RECT  7.225 2.730 7.455 3.455 ;
        RECT  6.290 2.730 7.225 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 -0.235 14.560 0.235 ;
        RECT  14.095 -0.235 14.325 1.245 ;
        RECT  12.940 -0.235 14.095 0.235 ;
        RECT  12.600 -0.235 12.940 1.180 ;
        RECT  11.460 -0.235 12.600 0.235 ;
        RECT  11.120 -0.235 11.460 0.465 ;
        RECT  9.530 -0.235 11.120 0.235 ;
        RECT  9.190 -0.235 9.530 0.465 ;
        RECT  5.570 -0.235 9.190 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  2.560 -0.235 5.230 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 3.685 14.560 4.155 ;
        RECT  14.095 2.255 14.325 4.155 ;
        RECT  12.940 3.685 14.095 4.155 ;
        RECT  12.600 3.250 12.940 4.155 ;
        RECT  11.345 3.685 12.600 4.155 ;
        RECT  11.005 3.250 11.345 4.155 ;
        RECT  9.745 3.685 11.005 4.155 ;
        RECT  9.405 3.190 9.745 4.155 ;
        RECT  6.995 3.685 9.405 4.155 ;
        RECT  6.655 3.190 6.995 4.155 ;
        RECT  2.385 3.685 6.655 4.155 ;
        RECT  2.045 3.455 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.895 1.600 13.125 3.020 ;
        RECT  11.120 2.790 12.895 3.020 ;
        RECT  11.410 0.695 11.640 1.940 ;
        RECT  8.715 0.695 11.410 0.925 ;
        RECT  10.890 1.155 11.120 3.020 ;
        RECT  9.675 1.155 10.890 1.385 ;
        RECT  10.465 2.540 10.890 2.770 ;
        RECT  10.360 1.670 10.590 2.260 ;
        RECT  10.235 2.540 10.465 3.370 ;
        RECT  9.695 2.030 10.360 2.260 ;
        RECT  9.465 2.030 9.695 2.960 ;
        RECT  9.445 1.155 9.675 1.750 ;
        RECT  7.915 2.730 9.465 2.960 ;
        RECT  8.945 1.520 9.445 1.750 ;
        RECT  8.715 2.270 8.910 2.500 ;
        RECT  8.485 0.465 8.715 2.500 ;
        RECT  7.435 0.990 8.485 1.220 ;
        RECT  7.685 1.615 7.915 2.960 ;
        RECT  7.140 1.615 7.685 1.845 ;
        RECT  6.910 0.985 7.140 1.845 ;
        RECT  6.505 2.270 7.060 2.500 ;
        RECT  6.715 0.985 6.910 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.075 2.460 5.735 2.690 ;
        RECT  3.845 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  3.140 0.465 4.145 0.695 ;
        RECT  1.650 2.980 3.935 3.210 ;
        RECT  3.615 0.990 3.845 2.690 ;
        RECT  3.490 0.990 3.615 1.220 ;
        RECT  3.320 2.460 3.615 2.690 ;
        RECT  2.910 0.465 3.140 1.205 ;
        RECT  2.095 0.975 2.910 1.205 ;
        RECT  1.865 0.975 2.095 2.680 ;
        RECT  1.520 0.975 1.865 1.205 ;
        RECT  1.520 2.450 1.865 2.680 ;
        RECT  1.310 2.980 1.650 3.455 ;
        RECT  0.465 2.980 1.310 3.210 ;
        RECT  0.345 0.975 0.530 1.205 ;
        RECT  0.345 2.470 0.465 3.210 ;
        RECT  0.235 0.975 0.345 3.210 ;
        RECT  0.115 0.975 0.235 2.810 ;
    END
END DFCND2BWP7T

MACRO DFCNQD1BWP7T
    CLASS CORE ;
    FOREIGN DFCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.850 0.470 12.180 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4158 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.725 3.385 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.700 1.540 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.455 3.225 8.570 3.455 ;
        RECT  7.225 2.730 7.455 3.455 ;
        RECT  6.290 2.730 7.225 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.365 -0.235 12.320 0.235 ;
        RECT  11.135 -0.235 11.365 1.290 ;
        RECT  8.875 -0.235 11.135 0.235 ;
        RECT  8.535 -0.235 8.875 0.465 ;
        RECT  5.570 -0.235 8.535 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  2.560 -0.235 5.230 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.330 3.685 12.320 4.155 ;
        RECT  11.100 2.255 11.330 4.155 ;
        RECT  9.705 3.685 11.100 4.155 ;
        RECT  9.365 3.190 9.705 4.155 ;
        RECT  6.995 3.685 9.365 4.155 ;
        RECT  6.655 3.190 6.995 4.155 ;
        RECT  2.385 3.685 6.655 4.155 ;
        RECT  2.045 3.455 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.840 1.600 11.605 1.940 ;
        RECT  10.620 0.990 10.840 2.795 ;
        RECT  10.610 0.465 10.620 2.795 ;
        RECT  10.390 0.465 10.610 1.220 ;
        RECT  10.520 2.565 10.610 2.795 ;
        RECT  10.290 2.565 10.520 3.375 ;
        RECT  9.700 0.990 10.390 1.220 ;
        RECT  10.150 1.565 10.380 2.330 ;
        RECT  9.655 2.100 10.150 2.330 ;
        RECT  9.470 0.990 9.700 1.845 ;
        RECT  9.425 2.100 9.655 2.960 ;
        RECT  8.825 1.615 9.470 1.845 ;
        RECT  7.915 2.730 9.425 2.960 ;
        RECT  8.495 0.990 8.815 1.220 ;
        RECT  8.495 2.270 8.815 2.500 ;
        RECT  8.265 0.990 8.495 2.500 ;
        RECT  7.535 0.990 8.265 1.220 ;
        RECT  7.685 1.615 7.915 2.960 ;
        RECT  7.140 1.615 7.685 1.845 ;
        RECT  6.910 0.985 7.140 1.845 ;
        RECT  6.505 2.270 7.060 2.500 ;
        RECT  6.750 0.985 6.910 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.075 2.460 5.735 2.690 ;
        RECT  3.845 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  3.140 0.465 4.145 0.695 ;
        RECT  1.650 2.980 3.935 3.210 ;
        RECT  3.615 0.990 3.845 2.690 ;
        RECT  3.490 0.990 3.615 1.220 ;
        RECT  3.320 2.460 3.615 2.690 ;
        RECT  2.910 0.465 3.140 1.205 ;
        RECT  2.095 0.975 2.910 1.205 ;
        RECT  1.865 0.975 2.095 2.680 ;
        RECT  1.520 0.975 1.865 1.205 ;
        RECT  1.520 2.450 1.865 2.680 ;
        RECT  1.310 2.980 1.650 3.455 ;
        RECT  0.465 2.980 1.310 3.210 ;
        RECT  0.345 0.975 0.530 1.205 ;
        RECT  0.345 2.470 0.465 3.210 ;
        RECT  0.235 0.975 0.345 3.210 ;
        RECT  0.115 0.975 0.235 2.810 ;
    END
END DFCNQD1BWP7T

MACRO DFCNQD2BWP7T
    CLASS CORE ;
    FOREIGN DFCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.925 1.065 12.180 2.730 ;
        RECT  11.900 0.470 11.925 3.310 ;
        RECT  11.690 0.470 11.900 1.295 ;
        RECT  11.695 2.500 11.900 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4158 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.725 3.385 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.700 1.540 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.500 3.225 8.965 3.455 ;
        RECT  7.270 2.730 7.500 3.455 ;
        RECT  6.290 2.730 7.270 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 -0.235 12.880 0.235 ;
        RECT  12.415 -0.235 12.645 1.235 ;
        RECT  11.260 -0.235 12.415 0.235 ;
        RECT  10.920 -0.235 11.260 0.755 ;
        RECT  8.825 -0.235 10.920 0.235 ;
        RECT  8.485 -0.235 8.825 0.465 ;
        RECT  5.570 -0.235 8.485 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  2.560 -0.235 5.230 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 3.685 12.880 4.155 ;
        RECT  12.415 2.255 12.645 4.155 ;
        RECT  11.255 3.685 12.415 4.155 ;
        RECT  10.915 3.090 11.255 4.155 ;
        RECT  9.715 3.685 10.915 4.155 ;
        RECT  9.375 3.190 9.715 4.155 ;
        RECT  7.040 3.685 9.375 4.155 ;
        RECT  6.700 3.190 7.040 4.155 ;
        RECT  2.385 3.685 6.700 4.155 ;
        RECT  2.045 3.455 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.190 1.600 11.590 1.940 ;
        RECT  10.960 0.990 11.190 2.795 ;
        RECT  10.505 0.990 10.960 1.220 ;
        RECT  10.475 2.565 10.960 2.795 ;
        RECT  10.275 0.465 10.505 1.220 ;
        RECT  10.275 1.565 10.505 2.260 ;
        RECT  10.245 2.565 10.475 3.375 ;
        RECT  9.645 0.990 10.275 1.220 ;
        RECT  9.655 2.030 10.275 2.260 ;
        RECT  9.425 2.030 9.655 2.960 ;
        RECT  9.415 0.990 9.645 1.760 ;
        RECT  7.960 2.730 9.425 2.960 ;
        RECT  8.870 1.530 9.415 1.760 ;
        RECT  8.535 0.990 8.810 1.220 ;
        RECT  8.535 2.270 8.790 2.500 ;
        RECT  8.305 0.990 8.535 2.500 ;
        RECT  7.480 0.990 8.305 1.220 ;
        RECT  7.730 1.670 7.960 2.960 ;
        RECT  7.185 1.670 7.730 1.900 ;
        RECT  6.955 0.985 7.185 1.900 ;
        RECT  6.505 2.270 7.105 2.500 ;
        RECT  6.715 0.985 6.955 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.075 2.460 5.735 2.690 ;
        RECT  3.845 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  3.140 0.465 4.145 0.695 ;
        RECT  1.650 2.980 3.935 3.210 ;
        RECT  3.615 0.990 3.845 2.690 ;
        RECT  3.490 0.990 3.615 1.220 ;
        RECT  3.320 2.460 3.615 2.690 ;
        RECT  2.910 0.465 3.140 1.205 ;
        RECT  2.095 0.975 2.910 1.205 ;
        RECT  1.865 0.975 2.095 2.680 ;
        RECT  1.520 0.975 1.865 1.205 ;
        RECT  1.520 2.450 1.865 2.680 ;
        RECT  1.310 2.980 1.650 3.455 ;
        RECT  0.465 2.980 1.310 3.210 ;
        RECT  0.345 0.975 0.530 1.205 ;
        RECT  0.345 2.470 0.465 3.210 ;
        RECT  0.235 0.975 0.345 3.210 ;
        RECT  0.115 0.975 0.235 2.810 ;
    END
END DFCNQD2BWP7T

MACRO DFD0BWP7T
    CLASS CORE ;
    FOREIGN DFD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.075 9.940 2.560 ;
        RECT  9.525 1.075 9.660 1.305 ;
        RECT  9.240 2.330 9.660 2.560 ;
        RECT  9.295 0.510 9.525 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.730 0.515 11.060 2.720 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 1.715 3.460 2.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 -0.235 11.200 0.235 ;
        RECT  9.960 -0.235 10.300 0.810 ;
        RECT  7.165 -0.235 9.960 0.235 ;
        RECT  6.825 -0.235 7.165 0.465 ;
        RECT  5.145 -0.235 6.825 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  2.560 -0.235 4.805 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.240 3.685 11.200 4.155 ;
        RECT  9.900 3.315 10.240 4.155 ;
        RECT  8.155 3.685 9.900 4.155 ;
        RECT  7.815 3.250 8.155 4.155 ;
        RECT  5.155 3.685 7.815 4.155 ;
        RECT  4.795 3.190 5.155 4.155 ;
        RECT  2.590 3.685 4.795 4.155 ;
        RECT  2.250 2.800 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.255 1.600 10.485 3.020 ;
        RECT  9.005 2.790 10.255 3.020 ;
        RECT  7.625 0.465 9.055 0.695 ;
        RECT  8.820 1.020 9.005 3.020 ;
        RECT  8.775 1.020 8.820 3.380 ;
        RECT  8.085 1.020 8.775 1.250 ;
        RECT  8.590 2.790 8.775 3.380 ;
        RECT  8.315 1.565 8.545 2.310 ;
        RECT  8.085 2.080 8.315 2.310 ;
        RECT  7.855 1.020 8.085 1.830 ;
        RECT  7.855 2.080 8.085 2.995 ;
        RECT  7.370 1.600 7.855 1.830 ;
        RECT  6.570 2.765 7.855 2.995 ;
        RECT  7.395 0.465 7.625 1.220 ;
        RECT  7.135 2.300 7.405 2.530 ;
        RECT  7.135 0.990 7.395 1.220 ;
        RECT  6.905 0.990 7.135 2.530 ;
        RECT  5.860 3.225 7.115 3.455 ;
        RECT  6.340 0.910 6.570 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.565 2.270 5.855 2.500 ;
        RECT  4.540 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.415 ;
        RECT  4.050 2.185 5.075 2.415 ;
        RECT  4.580 0.960 4.810 1.890 ;
        RECT  4.310 2.730 4.540 3.280 ;
        RECT  3.140 3.050 4.310 3.280 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.820 0.990 4.050 2.695 ;
        RECT  3.520 0.990 3.820 1.220 ;
        RECT  3.485 2.465 3.820 2.695 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.910 2.340 3.140 3.280 ;
        RECT  2.020 0.975 2.930 1.205 ;
        RECT  2.020 2.340 2.910 2.570 ;
        RECT  1.790 0.975 2.020 2.755 ;
        RECT  1.520 0.975 1.790 1.205 ;
        RECT  1.520 2.525 1.790 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.995 0.530 1.225 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.995 0.345 3.215 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFD0BWP7T

MACRO DFD1BWP7T
    CLASS CORE ;
    FOREIGN DFD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.075 9.940 2.560 ;
        RECT  9.525 1.075 9.660 1.305 ;
        RECT  9.240 2.330 9.660 2.560 ;
        RECT  9.295 0.480 9.525 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.730 0.470 11.060 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 1.715 3.460 2.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 -0.235 11.200 0.235 ;
        RECT  9.960 -0.235 10.300 0.810 ;
        RECT  7.165 -0.235 9.960 0.235 ;
        RECT  6.825 -0.235 7.165 0.465 ;
        RECT  5.145 -0.235 6.825 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  2.560 -0.235 4.805 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 3.685 11.200 4.155 ;
        RECT  9.960 3.250 10.300 4.155 ;
        RECT  8.155 3.685 9.960 4.155 ;
        RECT  7.815 3.250 8.155 4.155 ;
        RECT  5.155 3.685 7.815 4.155 ;
        RECT  4.795 3.190 5.155 4.155 ;
        RECT  2.590 3.685 4.795 4.155 ;
        RECT  2.250 2.800 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.255 1.600 10.485 3.020 ;
        RECT  9.005 2.790 10.255 3.020 ;
        RECT  7.625 0.465 9.055 0.695 ;
        RECT  8.820 1.020 9.005 3.020 ;
        RECT  8.775 1.020 8.820 3.380 ;
        RECT  8.085 1.020 8.775 1.250 ;
        RECT  8.590 2.565 8.775 3.380 ;
        RECT  8.315 1.565 8.545 2.310 ;
        RECT  8.085 2.080 8.315 2.310 ;
        RECT  7.855 1.020 8.085 1.830 ;
        RECT  7.855 2.080 8.085 2.995 ;
        RECT  7.370 1.600 7.855 1.830 ;
        RECT  6.570 2.765 7.855 2.995 ;
        RECT  7.395 0.465 7.625 1.220 ;
        RECT  7.135 2.300 7.405 2.530 ;
        RECT  7.135 0.990 7.395 1.220 ;
        RECT  6.905 0.990 7.135 2.530 ;
        RECT  5.860 3.225 7.115 3.455 ;
        RECT  6.340 0.910 6.570 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.565 2.270 5.855 2.500 ;
        RECT  4.540 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.415 ;
        RECT  4.050 2.185 5.075 2.415 ;
        RECT  4.580 0.960 4.810 1.890 ;
        RECT  4.310 2.730 4.540 3.280 ;
        RECT  3.140 3.050 4.310 3.280 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.820 0.990 4.050 2.695 ;
        RECT  3.520 0.990 3.820 1.220 ;
        RECT  3.485 2.465 3.820 2.695 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.910 2.340 3.140 3.280 ;
        RECT  2.020 0.975 2.930 1.205 ;
        RECT  2.020 2.340 2.910 2.570 ;
        RECT  1.790 0.975 2.020 2.755 ;
        RECT  1.520 0.975 1.790 1.205 ;
        RECT  1.520 2.525 1.790 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.995 0.530 1.225 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.995 0.345 3.215 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFD1BWP7T

MACRO DFD2BWP7T
    CLASS CORE ;
    FOREIGN DFD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.3211 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.200 0.465 10.545 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.925 1.055 12.180 2.690 ;
        RECT  11.900 0.465 11.925 3.310 ;
        RECT  11.690 0.465 11.900 1.285 ;
        RECT  11.695 2.460 11.900 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.715 3.445 2.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 -0.235 12.880 0.235 ;
        RECT  12.415 -0.235 12.645 1.245 ;
        RECT  11.260 -0.235 12.415 0.235 ;
        RECT  10.920 -0.235 11.260 1.180 ;
        RECT  9.780 -0.235 10.920 0.235 ;
        RECT  9.440 -0.235 9.780 0.465 ;
        RECT  8.150 -0.235 9.440 0.235 ;
        RECT  7.810 -0.235 8.150 0.465 ;
        RECT  5.130 -0.235 7.810 0.235 ;
        RECT  4.790 -0.235 5.130 0.730 ;
        RECT  2.560 -0.235 4.790 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 3.685 12.880 4.155 ;
        RECT  12.415 2.255 12.645 4.155 ;
        RECT  11.260 3.685 12.415 4.155 ;
        RECT  10.920 3.250 11.260 4.155 ;
        RECT  9.780 3.685 10.920 4.155 ;
        RECT  9.440 3.250 9.780 4.155 ;
        RECT  8.150 3.685 9.440 4.155 ;
        RECT  7.810 3.250 8.150 4.155 ;
        RECT  5.140 3.685 7.810 4.155 ;
        RECT  4.780 3.190 5.140 4.155 ;
        RECT  2.575 3.685 4.780 4.155 ;
        RECT  2.235 2.800 2.575 4.155 ;
        RECT  1.080 3.685 2.235 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.215 1.605 11.445 3.010 ;
        RECT  9.350 2.780 11.215 3.010 ;
        RECT  9.730 0.695 9.960 1.945 ;
        RECT  7.630 0.695 9.730 0.925 ;
        RECT  9.120 1.155 9.350 3.010 ;
        RECT  8.220 1.155 9.120 1.385 ;
        RECT  8.925 2.565 9.120 3.010 ;
        RECT  8.695 2.565 8.925 3.380 ;
        RECT  8.585 1.675 8.815 2.310 ;
        RECT  8.170 2.080 8.585 2.310 ;
        RECT  7.990 1.155 8.220 1.830 ;
        RECT  7.940 2.080 8.170 2.995 ;
        RECT  7.365 1.600 7.990 1.830 ;
        RECT  6.560 2.765 7.940 2.995 ;
        RECT  7.400 0.695 7.630 1.220 ;
        RECT  7.100 0.990 7.400 1.220 ;
        RECT  7.100 2.300 7.390 2.530 ;
        RECT  6.870 0.990 7.100 2.530 ;
        RECT  5.845 3.225 7.005 3.455 ;
        RECT  6.325 0.910 6.560 2.995 ;
        RECT  5.840 0.960 6.070 2.500 ;
        RECT  5.615 2.730 5.845 3.455 ;
        RECT  4.795 0.960 5.840 1.190 ;
        RECT  5.550 2.270 5.840 2.500 ;
        RECT  4.525 2.730 5.615 2.960 ;
        RECT  5.290 1.560 5.595 1.900 ;
        RECT  5.060 1.560 5.290 2.415 ;
        RECT  4.035 2.185 5.060 2.415 ;
        RECT  4.565 0.960 4.795 1.890 ;
        RECT  4.295 2.730 4.525 3.280 ;
        RECT  3.125 3.050 4.295 3.280 ;
        RECT  3.145 0.465 4.115 0.695 ;
        RECT  3.805 0.990 4.035 2.695 ;
        RECT  3.505 0.990 3.805 1.220 ;
        RECT  3.470 2.465 3.805 2.695 ;
        RECT  2.915 0.465 3.145 1.205 ;
        RECT  2.895 2.340 3.125 3.280 ;
        RECT  2.000 0.975 2.915 1.205 ;
        RECT  2.000 2.340 2.895 2.570 ;
        RECT  1.770 0.975 2.000 2.755 ;
        RECT  1.520 0.975 1.770 1.205 ;
        RECT  1.520 2.525 1.770 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.995 0.530 1.225 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.995 0.345 3.215 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFD2BWP7T

MACRO DFKCND0BWP7T
    CLASS CORE ;
    FOREIGN DFKCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.780 1.075 11.060 2.560 ;
        RECT  10.645 1.075 10.780 1.305 ;
        RECT  10.360 2.330 10.780 2.560 ;
        RECT  10.415 0.510 10.645 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.850 0.515 12.180 2.715 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.735 3.855 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.760 0.980 2.710 ;
        RECT  0.590 1.760 0.700 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2502 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.735 2.675 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.420 -0.235 12.320 0.235 ;
        RECT  11.080 -0.235 11.420 0.810 ;
        RECT  8.285 -0.235 11.080 0.235 ;
        RECT  7.945 -0.235 8.285 0.465 ;
        RECT  6.265 -0.235 7.945 0.235 ;
        RECT  5.925 -0.235 6.265 0.730 ;
        RECT  2.800 -0.235 5.925 0.235 ;
        RECT  2.460 -0.235 2.800 0.730 ;
        RECT  1.285 -0.235 2.460 0.235 ;
        RECT  0.945 -0.235 1.285 0.745 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.380 3.685 12.320 4.155 ;
        RECT  11.040 3.335 11.380 4.155 ;
        RECT  9.275 3.685 11.040 4.155 ;
        RECT  8.935 3.250 9.275 4.155 ;
        RECT  6.265 3.685 8.935 4.155 ;
        RECT  5.925 3.190 6.265 4.155 ;
        RECT  3.300 3.685 5.925 4.155 ;
        RECT  2.960 2.885 3.300 4.155 ;
        RECT  1.080 3.685 2.960 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.375 1.600 11.605 3.020 ;
        RECT  10.125 2.790 11.375 3.020 ;
        RECT  8.745 0.465 10.170 0.695 ;
        RECT  9.940 0.990 10.125 3.020 ;
        RECT  9.895 0.990 9.940 3.380 ;
        RECT  9.205 0.990 9.895 1.220 ;
        RECT  9.710 2.790 9.895 3.380 ;
        RECT  9.435 1.565 9.665 2.310 ;
        RECT  9.205 2.080 9.435 2.310 ;
        RECT  8.975 0.990 9.205 1.830 ;
        RECT  8.975 2.080 9.205 2.995 ;
        RECT  8.490 1.600 8.975 1.830 ;
        RECT  7.690 2.765 8.975 2.995 ;
        RECT  8.515 0.465 8.745 1.220 ;
        RECT  8.255 2.300 8.525 2.530 ;
        RECT  8.255 0.990 8.515 1.220 ;
        RECT  8.025 0.990 8.255 2.530 ;
        RECT  6.980 3.225 8.235 3.455 ;
        RECT  7.460 0.910 7.690 2.995 ;
        RECT  6.980 0.960 7.210 2.500 ;
        RECT  5.960 0.960 6.980 1.190 ;
        RECT  6.685 2.270 6.980 2.500 ;
        RECT  6.750 2.730 6.980 3.455 ;
        RECT  5.560 2.730 6.750 2.960 ;
        RECT  6.455 1.560 6.730 1.900 ;
        RECT  6.225 1.560 6.455 2.415 ;
        RECT  4.980 2.185 6.225 2.415 ;
        RECT  5.730 0.960 5.960 1.890 ;
        RECT  5.330 2.730 5.560 3.345 ;
        RECT  4.520 3.115 5.330 3.345 ;
        RECT  4.520 0.465 5.280 0.700 ;
        RECT  4.750 0.935 4.980 2.750 ;
        RECT  4.290 0.465 4.520 3.345 ;
        RECT  1.520 0.980 4.290 1.210 ;
        RECT  2.200 2.410 4.060 2.640 ;
        RECT  1.520 2.440 1.840 2.670 ;
        RECT  1.330 2.995 1.675 3.455 ;
        RECT  1.290 0.980 1.520 2.670 ;
        RECT  0.465 2.995 1.330 3.225 ;
        RECT  0.360 0.975 0.520 1.205 ;
        RECT  0.360 2.505 0.465 3.225 ;
        RECT  0.235 0.975 0.360 3.225 ;
        RECT  0.130 0.975 0.235 2.790 ;
    END
END DFKCND0BWP7T

MACRO DFKCND1BWP7T
    CLASS CORE ;
    FOREIGN DFKCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.780 1.075 11.060 2.560 ;
        RECT  10.645 1.075 10.780 1.305 ;
        RECT  10.360 2.330 10.780 2.560 ;
        RECT  10.415 0.480 10.645 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.850 0.470 12.180 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.735 3.855 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.760 0.980 2.710 ;
        RECT  0.590 1.760 0.700 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2502 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.735 2.675 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.420 -0.235 12.320 0.235 ;
        RECT  11.080 -0.235 11.420 0.810 ;
        RECT  8.285 -0.235 11.080 0.235 ;
        RECT  7.945 -0.235 8.285 0.465 ;
        RECT  6.265 -0.235 7.945 0.235 ;
        RECT  5.925 -0.235 6.265 0.730 ;
        RECT  2.800 -0.235 5.925 0.235 ;
        RECT  2.460 -0.235 2.800 0.730 ;
        RECT  1.285 -0.235 2.460 0.235 ;
        RECT  0.945 -0.235 1.285 0.745 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.420 3.685 12.320 4.155 ;
        RECT  11.080 3.250 11.420 4.155 ;
        RECT  9.275 3.685 11.080 4.155 ;
        RECT  8.935 3.250 9.275 4.155 ;
        RECT  6.265 3.685 8.935 4.155 ;
        RECT  5.925 3.190 6.265 4.155 ;
        RECT  3.300 3.685 5.925 4.155 ;
        RECT  2.960 2.885 3.300 4.155 ;
        RECT  1.080 3.685 2.960 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.375 1.600 11.605 3.020 ;
        RECT  10.125 2.790 11.375 3.020 ;
        RECT  8.745 0.465 10.170 0.695 ;
        RECT  9.940 1.020 10.125 3.020 ;
        RECT  9.895 1.020 9.940 3.380 ;
        RECT  9.205 1.020 9.895 1.250 ;
        RECT  9.710 2.565 9.895 3.380 ;
        RECT  9.435 1.565 9.665 2.310 ;
        RECT  9.205 2.080 9.435 2.310 ;
        RECT  8.975 1.020 9.205 1.830 ;
        RECT  8.975 2.080 9.205 2.995 ;
        RECT  8.490 1.600 8.975 1.830 ;
        RECT  7.690 2.765 8.975 2.995 ;
        RECT  8.515 0.465 8.745 1.220 ;
        RECT  8.255 2.300 8.525 2.530 ;
        RECT  8.255 0.990 8.515 1.220 ;
        RECT  8.025 0.990 8.255 2.530 ;
        RECT  6.980 3.225 8.235 3.455 ;
        RECT  7.460 0.910 7.690 2.995 ;
        RECT  6.980 0.960 7.210 2.500 ;
        RECT  5.960 0.960 6.980 1.190 ;
        RECT  6.685 2.270 6.980 2.500 ;
        RECT  6.750 2.730 6.980 3.455 ;
        RECT  5.560 2.730 6.750 2.960 ;
        RECT  6.455 1.560 6.730 1.900 ;
        RECT  6.225 1.560 6.455 2.415 ;
        RECT  4.980 2.185 6.225 2.415 ;
        RECT  5.730 0.960 5.960 1.890 ;
        RECT  5.330 2.730 5.560 3.345 ;
        RECT  4.520 3.115 5.330 3.345 ;
        RECT  4.520 0.465 5.280 0.700 ;
        RECT  4.750 0.935 4.980 2.750 ;
        RECT  4.290 0.465 4.520 3.345 ;
        RECT  1.520 0.980 4.290 1.210 ;
        RECT  2.200 2.410 4.060 2.640 ;
        RECT  1.520 2.440 1.840 2.670 ;
        RECT  1.330 2.995 1.675 3.455 ;
        RECT  1.290 0.980 1.520 2.670 ;
        RECT  0.465 2.995 1.330 3.225 ;
        RECT  0.360 0.975 0.520 1.205 ;
        RECT  0.360 2.505 0.465 3.225 ;
        RECT  0.235 0.975 0.360 3.225 ;
        RECT  0.130 0.975 0.235 2.790 ;
    END
END DFKCND1BWP7T

MACRO DFKCND2BWP7T
    CLASS CORE ;
    FOREIGN DFKCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.320 0.465 11.665 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.045 1.055 13.300 2.690 ;
        RECT  13.020 0.465 13.045 3.310 ;
        RECT  12.810 0.465 13.020 1.285 ;
        RECT  12.815 2.460 13.020 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.735 3.855 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.760 0.980 2.710 ;
        RECT  0.590 1.760 0.700 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2502 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.735 2.675 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.765 -0.235 14.000 0.235 ;
        RECT  13.535 -0.235 13.765 1.245 ;
        RECT  12.380 -0.235 13.535 0.235 ;
        RECT  12.040 -0.235 12.380 1.180 ;
        RECT  10.900 -0.235 12.040 0.235 ;
        RECT  10.560 -0.235 10.900 0.465 ;
        RECT  9.285 -0.235 10.560 0.235 ;
        RECT  8.945 -0.235 9.285 0.465 ;
        RECT  6.265 -0.235 8.945 0.235 ;
        RECT  5.925 -0.235 6.265 0.730 ;
        RECT  2.800 -0.235 5.925 0.235 ;
        RECT  2.460 -0.235 2.800 0.730 ;
        RECT  1.285 -0.235 2.460 0.235 ;
        RECT  0.945 -0.235 1.285 0.745 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.765 3.685 14.000 4.155 ;
        RECT  13.535 2.255 13.765 4.155 ;
        RECT  12.380 3.685 13.535 4.155 ;
        RECT  12.040 3.250 12.380 4.155 ;
        RECT  10.900 3.685 12.040 4.155 ;
        RECT  10.560 3.250 10.900 4.155 ;
        RECT  9.285 3.685 10.560 4.155 ;
        RECT  8.945 3.250 9.285 4.155 ;
        RECT  6.265 3.685 8.945 4.155 ;
        RECT  5.925 3.190 6.265 4.155 ;
        RECT  3.300 3.685 5.925 4.155 ;
        RECT  2.960 2.885 3.300 4.155 ;
        RECT  1.080 3.685 2.960 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.335 1.605 12.565 3.010 ;
        RECT  10.485 2.780 12.335 3.010 ;
        RECT  10.850 0.695 11.080 1.945 ;
        RECT  8.765 0.695 10.850 0.925 ;
        RECT  10.255 1.155 10.485 3.010 ;
        RECT  9.355 1.155 10.255 1.385 ;
        RECT  10.060 2.565 10.255 3.010 ;
        RECT  9.830 2.565 10.060 3.380 ;
        RECT  9.720 1.675 9.950 2.310 ;
        RECT  9.305 2.080 9.720 2.310 ;
        RECT  9.125 1.155 9.355 1.830 ;
        RECT  9.075 2.080 9.305 2.995 ;
        RECT  8.500 1.600 9.125 1.830 ;
        RECT  7.695 2.765 9.075 2.995 ;
        RECT  8.535 0.695 8.765 1.220 ;
        RECT  8.235 0.990 8.535 1.220 ;
        RECT  8.235 2.300 8.525 2.530 ;
        RECT  8.005 0.990 8.235 2.530 ;
        RECT  6.980 3.225 8.140 3.455 ;
        RECT  7.460 0.910 7.695 2.995 ;
        RECT  6.980 0.960 7.210 2.500 ;
        RECT  5.960 0.960 6.980 1.190 ;
        RECT  6.685 2.270 6.980 2.500 ;
        RECT  6.750 2.730 6.980 3.455 ;
        RECT  5.560 2.730 6.750 2.960 ;
        RECT  6.455 1.560 6.730 1.900 ;
        RECT  6.225 1.560 6.455 2.415 ;
        RECT  4.980 2.185 6.225 2.415 ;
        RECT  5.730 0.960 5.960 1.890 ;
        RECT  5.330 2.730 5.560 3.345 ;
        RECT  4.520 3.115 5.330 3.345 ;
        RECT  4.520 0.465 5.280 0.700 ;
        RECT  4.750 0.935 4.980 2.750 ;
        RECT  4.290 0.465 4.520 3.345 ;
        RECT  1.520 0.980 4.290 1.210 ;
        RECT  2.200 2.410 4.060 2.640 ;
        RECT  1.520 2.440 1.840 2.670 ;
        RECT  1.330 2.995 1.675 3.455 ;
        RECT  1.290 0.980 1.520 2.670 ;
        RECT  0.465 2.995 1.330 3.225 ;
        RECT  0.360 0.975 0.520 1.205 ;
        RECT  0.360 2.505 0.465 3.225 ;
        RECT  0.235 0.975 0.360 3.225 ;
        RECT  0.130 0.975 0.235 2.790 ;
    END
END DFKCND2BWP7T

MACRO DFKCNQD1BWP7T
    CLASS CORE ;
    FOREIGN DFKCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.730 0.470 11.060 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.735 3.855 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.760 0.980 2.710 ;
        RECT  0.590 1.760 0.700 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2502 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.735 2.675 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 -0.235 11.200 0.235 ;
        RECT  9.960 -0.235 10.300 0.765 ;
        RECT  8.285 -0.235 9.960 0.235 ;
        RECT  7.945 -0.235 8.285 0.465 ;
        RECT  6.245 -0.235 7.945 0.235 ;
        RECT  5.905 -0.235 6.245 0.730 ;
        RECT  2.800 -0.235 5.905 0.235 ;
        RECT  2.460 -0.235 2.800 0.730 ;
        RECT  1.285 -0.235 2.460 0.235 ;
        RECT  0.945 -0.235 1.285 0.745 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 3.685 11.200 4.155 ;
        RECT  9.960 3.250 10.300 4.155 ;
        RECT  9.040 3.685 9.960 4.155 ;
        RECT  8.700 2.590 9.040 4.155 ;
        RECT  6.245 3.685 8.700 4.155 ;
        RECT  5.905 3.190 6.245 4.155 ;
        RECT  3.300 3.685 5.905 4.155 ;
        RECT  2.960 2.885 3.300 4.155 ;
        RECT  1.080 3.685 2.960 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.205 1.020 10.435 2.755 ;
        RECT  9.545 1.020 10.205 1.250 ;
        RECT  9.415 2.525 10.205 2.755 ;
        RECT  9.315 0.495 9.545 1.250 ;
        RECT  9.100 1.565 9.330 2.310 ;
        RECT  8.655 1.020 9.315 1.250 ;
        RECT  7.670 2.080 9.100 2.310 ;
        RECT  8.315 1.020 8.655 1.830 ;
        RECT  6.960 3.225 8.100 3.455 ;
        RECT  7.440 0.910 7.670 2.850 ;
        RECT  6.960 0.960 7.190 2.500 ;
        RECT  5.940 0.960 6.960 1.190 ;
        RECT  6.665 2.270 6.960 2.500 ;
        RECT  6.730 2.730 6.960 3.455 ;
        RECT  5.540 2.730 6.730 2.960 ;
        RECT  6.435 1.560 6.710 1.900 ;
        RECT  6.205 1.560 6.435 2.415 ;
        RECT  4.960 2.185 6.205 2.415 ;
        RECT  5.710 0.960 5.940 1.890 ;
        RECT  5.310 2.730 5.540 3.345 ;
        RECT  4.500 3.115 5.310 3.345 ;
        RECT  4.500 0.465 5.260 0.700 ;
        RECT  4.730 0.935 4.960 2.750 ;
        RECT  4.270 0.465 4.500 3.345 ;
        RECT  1.520 0.980 4.270 1.210 ;
        RECT  3.775 2.410 4.005 2.750 ;
        RECT  2.200 2.410 3.775 2.640 ;
        RECT  1.520 2.440 1.840 2.670 ;
        RECT  1.330 2.995 1.675 3.455 ;
        RECT  1.290 0.980 1.520 2.670 ;
        RECT  0.465 2.995 1.330 3.225 ;
        RECT  0.360 0.975 0.520 1.205 ;
        RECT  0.360 2.505 0.465 3.225 ;
        RECT  0.235 0.975 0.360 3.225 ;
        RECT  0.130 0.975 0.235 2.790 ;
    END
END DFKCNQD1BWP7T

MACRO DFKCNQD2BWP7T
    CLASS CORE ;
    FOREIGN DFKCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.805 1.055 11.060 2.730 ;
        RECT  10.780 0.470 10.805 3.310 ;
        RECT  10.575 0.470 10.780 1.290 ;
        RECT  10.570 2.500 10.780 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.735 3.785 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.760 0.980 2.710 ;
        RECT  0.590 1.760 0.700 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2502 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.735 2.675 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.525 -0.235 11.760 0.235 ;
        RECT  11.295 -0.235 11.525 1.255 ;
        RECT  10.140 -0.235 11.295 0.235 ;
        RECT  9.800 -0.235 10.140 0.765 ;
        RECT  8.125 -0.235 9.800 0.235 ;
        RECT  7.785 -0.235 8.125 0.465 ;
        RECT  6.085 -0.235 7.785 0.235 ;
        RECT  5.745 -0.235 6.085 0.730 ;
        RECT  2.750 -0.235 5.745 0.235 ;
        RECT  2.410 -0.235 2.750 0.730 ;
        RECT  1.285 -0.235 2.410 0.235 ;
        RECT  0.945 -0.235 1.285 0.745 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.525 3.685 11.760 4.155 ;
        RECT  11.295 2.255 11.525 4.155 ;
        RECT  10.140 3.685 11.295 4.155 ;
        RECT  9.800 3.250 10.140 4.155 ;
        RECT  8.880 3.685 9.800 4.155 ;
        RECT  8.540 2.590 8.880 4.155 ;
        RECT  6.085 3.685 8.540 4.155 ;
        RECT  5.745 3.190 6.085 4.155 ;
        RECT  3.110 3.685 5.745 4.155 ;
        RECT  2.770 3.170 3.110 4.155 ;
        RECT  1.080 3.685 2.770 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.045 1.020 10.275 2.755 ;
        RECT  9.385 1.020 10.045 1.250 ;
        RECT  9.255 2.525 10.045 2.755 ;
        RECT  9.155 0.495 9.385 1.250 ;
        RECT  8.940 1.565 9.170 2.310 ;
        RECT  8.495 1.020 9.155 1.250 ;
        RECT  7.510 2.080 8.940 2.310 ;
        RECT  8.155 1.020 8.495 1.830 ;
        RECT  6.800 3.225 7.940 3.455 ;
        RECT  7.280 0.910 7.510 2.850 ;
        RECT  6.800 0.960 7.030 2.500 ;
        RECT  5.780 0.960 6.800 1.190 ;
        RECT  6.505 2.270 6.800 2.500 ;
        RECT  6.570 2.730 6.800 3.455 ;
        RECT  5.380 2.730 6.570 2.960 ;
        RECT  6.275 1.560 6.550 1.900 ;
        RECT  6.045 1.560 6.275 2.415 ;
        RECT  4.800 2.185 6.045 2.415 ;
        RECT  5.550 0.960 5.780 1.890 ;
        RECT  5.150 2.730 5.380 3.345 ;
        RECT  4.340 3.115 5.150 3.345 ;
        RECT  4.340 0.465 5.100 0.700 ;
        RECT  4.570 0.935 4.800 2.750 ;
        RECT  4.110 0.465 4.340 3.345 ;
        RECT  1.520 0.980 4.110 1.210 ;
        RECT  3.615 2.410 3.845 2.750 ;
        RECT  2.200 2.410 3.615 2.640 ;
        RECT  1.520 2.440 1.840 2.670 ;
        RECT  1.330 2.995 1.675 3.455 ;
        RECT  1.290 0.980 1.520 2.670 ;
        RECT  0.465 2.995 1.330 3.225 ;
        RECT  0.360 0.975 0.520 1.205 ;
        RECT  0.360 2.505 0.465 3.225 ;
        RECT  0.235 0.975 0.360 3.225 ;
        RECT  0.130 0.975 0.235 2.790 ;
    END
END DFKCNQD2BWP7T

MACRO DFKSND0BWP7T
    CLASS CORE ;
    FOREIGN DFKSND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.980 2.150 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.075 12.180 2.560 ;
        RECT  11.765 1.075 11.900 1.305 ;
        RECT  11.480 2.330 11.900 2.560 ;
        RECT  11.535 0.510 11.765 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.970 0.515 13.300 2.720 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 1.210 2.660 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 1.760 4.340 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 -0.235 13.440 0.235 ;
        RECT  12.200 -0.235 12.540 0.810 ;
        RECT  9.405 -0.235 12.200 0.235 ;
        RECT  9.065 -0.235 9.405 0.465 ;
        RECT  7.385 -0.235 9.065 0.235 ;
        RECT  7.045 -0.235 7.385 0.730 ;
        RECT  2.855 -0.235 7.045 0.235 ;
        RECT  2.515 -0.235 2.855 0.465 ;
        RECT  1.280 -0.235 2.515 0.235 ;
        RECT  0.940 -0.235 1.280 0.745 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.480 3.685 13.440 4.155 ;
        RECT  12.140 3.315 12.480 4.155 ;
        RECT  10.395 3.685 12.140 4.155 ;
        RECT  10.055 3.250 10.395 4.155 ;
        RECT  7.385 3.685 10.055 4.155 ;
        RECT  7.045 3.190 7.385 4.155 ;
        RECT  3.615 3.685 7.045 4.155 ;
        RECT  3.275 3.455 3.615 4.155 ;
        RECT  1.300 3.685 3.275 4.155 ;
        RECT  0.960 3.025 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.495 1.600 12.725 3.020 ;
        RECT  11.245 2.790 12.495 3.020 ;
        RECT  9.865 0.465 11.295 0.695 ;
        RECT  11.060 1.020 11.245 3.020 ;
        RECT  11.015 1.020 11.060 3.380 ;
        RECT  10.325 1.020 11.015 1.250 ;
        RECT  10.830 2.790 11.015 3.380 ;
        RECT  10.555 1.565 10.785 2.310 ;
        RECT  10.325 2.080 10.555 2.310 ;
        RECT  10.095 1.020 10.325 1.830 ;
        RECT  10.095 2.080 10.325 2.995 ;
        RECT  9.610 1.600 10.095 1.830 ;
        RECT  8.810 2.765 10.095 2.995 ;
        RECT  9.635 0.465 9.865 1.220 ;
        RECT  9.375 2.300 9.645 2.530 ;
        RECT  9.375 0.990 9.635 1.220 ;
        RECT  9.145 0.990 9.375 2.530 ;
        RECT  8.100 3.225 9.355 3.455 ;
        RECT  8.580 0.910 8.810 2.995 ;
        RECT  8.100 0.960 8.330 2.500 ;
        RECT  7.080 0.960 8.100 1.190 ;
        RECT  7.805 2.270 8.100 2.500 ;
        RECT  7.870 2.730 8.100 3.455 ;
        RECT  6.665 2.730 7.870 2.960 ;
        RECT  7.575 1.560 7.850 1.900 ;
        RECT  7.345 1.560 7.575 2.415 ;
        RECT  6.100 2.185 7.345 2.415 ;
        RECT  6.850 0.960 7.080 1.890 ;
        RECT  6.435 2.730 6.665 3.455 ;
        RECT  5.315 3.225 6.435 3.455 ;
        RECT  5.870 0.935 6.100 2.850 ;
        RECT  5.095 0.490 5.435 2.575 ;
        RECT  5.085 2.805 5.315 3.455 ;
        RECT  3.710 0.490 5.095 0.720 ;
        RECT  4.845 2.805 5.085 3.035 ;
        RECT  4.615 0.970 4.845 3.035 ;
        RECT  4.380 0.970 4.615 1.200 ;
        RECT  4.380 2.440 4.615 2.670 ;
        RECT  4.110 3.225 4.470 3.455 ;
        RECT  3.880 2.570 4.110 3.455 ;
        RECT  3.190 2.570 3.880 2.800 ;
        RECT  3.475 0.490 3.710 0.925 ;
        RECT  2.025 0.695 3.475 0.925 ;
        RECT  3.190 1.155 3.390 1.385 ;
        RECT  2.960 1.155 3.190 2.800 ;
        RECT  2.285 2.565 2.515 3.375 ;
        RECT  2.025 2.565 2.285 2.795 ;
        RECT  1.795 0.470 2.025 2.795 ;
        RECT  1.255 0.975 1.485 2.655 ;
        RECT  0.180 0.975 1.255 1.205 ;
        RECT  0.180 2.425 1.255 2.655 ;
    END
END DFKSND0BWP7T

MACRO DFKSND1BWP7T
    CLASS CORE ;
    FOREIGN DFKSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.980 2.150 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.075 12.180 2.560 ;
        RECT  11.765 1.075 11.900 1.305 ;
        RECT  11.480 2.330 11.900 2.560 ;
        RECT  11.535 0.480 11.765 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.970 0.470 13.300 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 1.210 2.660 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 1.760 4.340 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 -0.235 13.440 0.235 ;
        RECT  12.200 -0.235 12.540 0.810 ;
        RECT  9.405 -0.235 12.200 0.235 ;
        RECT  9.065 -0.235 9.405 0.465 ;
        RECT  7.385 -0.235 9.065 0.235 ;
        RECT  7.045 -0.235 7.385 0.730 ;
        RECT  2.855 -0.235 7.045 0.235 ;
        RECT  2.515 -0.235 2.855 0.465 ;
        RECT  1.280 -0.235 2.515 0.235 ;
        RECT  0.940 -0.235 1.280 0.745 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 3.685 13.440 4.155 ;
        RECT  12.200 3.250 12.540 4.155 ;
        RECT  10.395 3.685 12.200 4.155 ;
        RECT  10.055 3.250 10.395 4.155 ;
        RECT  7.385 3.685 10.055 4.155 ;
        RECT  7.045 3.190 7.385 4.155 ;
        RECT  3.615 3.685 7.045 4.155 ;
        RECT  3.275 3.455 3.615 4.155 ;
        RECT  1.300 3.685 3.275 4.155 ;
        RECT  0.960 3.025 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.495 1.600 12.725 3.020 ;
        RECT  11.245 2.790 12.495 3.020 ;
        RECT  9.865 0.465 11.290 0.695 ;
        RECT  11.060 0.990 11.245 3.020 ;
        RECT  11.015 0.990 11.060 3.380 ;
        RECT  10.325 0.990 11.015 1.220 ;
        RECT  10.830 2.565 11.015 3.380 ;
        RECT  10.555 1.565 10.785 2.310 ;
        RECT  10.325 2.080 10.555 2.310 ;
        RECT  10.095 0.990 10.325 1.850 ;
        RECT  10.095 2.080 10.325 2.995 ;
        RECT  9.610 1.620 10.095 1.850 ;
        RECT  8.810 2.765 10.095 2.995 ;
        RECT  9.635 0.465 9.865 1.220 ;
        RECT  9.375 2.300 9.645 2.530 ;
        RECT  9.375 0.990 9.635 1.220 ;
        RECT  9.145 0.990 9.375 2.530 ;
        RECT  8.100 3.225 9.355 3.455 ;
        RECT  8.580 0.935 8.810 2.995 ;
        RECT  8.100 0.960 8.330 2.500 ;
        RECT  7.080 0.960 8.100 1.190 ;
        RECT  7.805 2.270 8.100 2.500 ;
        RECT  7.870 2.730 8.100 3.455 ;
        RECT  6.665 2.730 7.870 2.960 ;
        RECT  7.575 1.560 7.850 1.900 ;
        RECT  7.345 1.560 7.575 2.415 ;
        RECT  6.100 2.185 7.345 2.415 ;
        RECT  6.850 0.960 7.080 1.890 ;
        RECT  6.435 2.730 6.665 3.455 ;
        RECT  5.315 3.225 6.435 3.455 ;
        RECT  5.870 0.935 6.100 2.850 ;
        RECT  5.095 0.490 5.435 2.575 ;
        RECT  5.085 2.805 5.315 3.455 ;
        RECT  3.710 0.490 5.095 0.720 ;
        RECT  4.845 2.805 5.085 3.035 ;
        RECT  4.615 0.970 4.845 3.035 ;
        RECT  4.380 0.970 4.615 1.200 ;
        RECT  4.380 2.440 4.615 2.670 ;
        RECT  4.110 3.225 4.470 3.455 ;
        RECT  3.880 2.570 4.110 3.455 ;
        RECT  3.190 2.570 3.880 2.800 ;
        RECT  3.475 0.490 3.710 0.925 ;
        RECT  2.025 0.695 3.475 0.925 ;
        RECT  3.190 1.155 3.390 1.385 ;
        RECT  2.960 1.155 3.190 2.800 ;
        RECT  2.285 2.565 2.515 3.375 ;
        RECT  2.025 2.565 2.285 2.795 ;
        RECT  1.795 0.470 2.025 2.795 ;
        RECT  1.255 0.975 1.485 2.655 ;
        RECT  0.180 0.975 1.255 1.205 ;
        RECT  0.180 2.425 1.255 2.655 ;
    END
END DFKSND1BWP7T

MACRO DFKSND2BWP7T
    CLASS CORE ;
    FOREIGN DFKSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.755 0.980 2.150 ;
        END
    END SN
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.440 0.465 12.785 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.165 1.055 14.420 2.690 ;
        RECT  14.140 0.465 14.165 3.310 ;
        RECT  13.930 0.465 14.140 1.285 ;
        RECT  13.935 2.460 14.140 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 1.210 2.660 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 1.760 4.340 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.885 -0.235 15.120 0.235 ;
        RECT  14.655 -0.235 14.885 1.245 ;
        RECT  13.500 -0.235 14.655 0.235 ;
        RECT  13.160 -0.235 13.500 1.180 ;
        RECT  12.020 -0.235 13.160 0.235 ;
        RECT  11.680 -0.235 12.020 0.465 ;
        RECT  10.405 -0.235 11.680 0.235 ;
        RECT  10.065 -0.235 10.405 0.465 ;
        RECT  7.385 -0.235 10.065 0.235 ;
        RECT  7.045 -0.235 7.385 0.730 ;
        RECT  2.855 -0.235 7.045 0.235 ;
        RECT  2.515 -0.235 2.855 0.465 ;
        RECT  1.280 -0.235 2.515 0.235 ;
        RECT  0.940 -0.235 1.280 0.745 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.885 3.685 15.120 4.155 ;
        RECT  14.655 2.255 14.885 4.155 ;
        RECT  13.500 3.685 14.655 4.155 ;
        RECT  13.160 3.250 13.500 4.155 ;
        RECT  12.020 3.685 13.160 4.155 ;
        RECT  11.680 3.250 12.020 4.155 ;
        RECT  10.405 3.685 11.680 4.155 ;
        RECT  10.065 3.250 10.405 4.155 ;
        RECT  7.385 3.685 10.065 4.155 ;
        RECT  7.045 3.190 7.385 4.155 ;
        RECT  3.615 3.685 7.045 4.155 ;
        RECT  3.275 3.455 3.615 4.155 ;
        RECT  1.300 3.685 3.275 4.155 ;
        RECT  0.960 3.025 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.455 1.605 13.685 3.010 ;
        RECT  11.605 2.780 13.455 3.010 ;
        RECT  11.970 0.695 12.200 1.945 ;
        RECT  9.885 0.695 11.970 0.925 ;
        RECT  11.375 1.155 11.605 3.010 ;
        RECT  10.475 1.155 11.375 1.385 ;
        RECT  11.180 2.565 11.375 3.010 ;
        RECT  10.950 2.565 11.180 3.380 ;
        RECT  10.840 1.675 11.070 2.310 ;
        RECT  10.425 2.080 10.840 2.310 ;
        RECT  10.245 1.155 10.475 1.830 ;
        RECT  10.195 2.080 10.425 2.995 ;
        RECT  9.620 1.600 10.245 1.830 ;
        RECT  8.815 2.765 10.195 2.995 ;
        RECT  9.655 0.695 9.885 1.220 ;
        RECT  9.355 0.990 9.655 1.220 ;
        RECT  9.355 2.300 9.645 2.530 ;
        RECT  9.125 0.990 9.355 2.530 ;
        RECT  8.100 3.225 9.260 3.455 ;
        RECT  8.580 0.910 8.815 2.995 ;
        RECT  8.100 0.960 8.330 2.500 ;
        RECT  7.080 0.960 8.100 1.190 ;
        RECT  7.805 2.270 8.100 2.500 ;
        RECT  7.870 2.730 8.100 3.455 ;
        RECT  6.665 2.730 7.870 2.960 ;
        RECT  7.575 1.560 7.850 1.900 ;
        RECT  7.345 1.560 7.575 2.415 ;
        RECT  6.100 2.185 7.345 2.415 ;
        RECT  6.850 0.960 7.080 1.890 ;
        RECT  6.435 2.730 6.665 3.455 ;
        RECT  5.315 3.225 6.435 3.455 ;
        RECT  5.870 0.935 6.100 2.850 ;
        RECT  5.095 0.490 5.435 2.575 ;
        RECT  5.085 2.805 5.315 3.455 ;
        RECT  3.710 0.490 5.095 0.720 ;
        RECT  4.845 2.805 5.085 3.035 ;
        RECT  4.615 0.970 4.845 3.035 ;
        RECT  4.380 0.970 4.615 1.200 ;
        RECT  4.380 2.440 4.615 2.670 ;
        RECT  4.110 3.225 4.470 3.455 ;
        RECT  3.880 2.570 4.110 3.455 ;
        RECT  3.190 2.570 3.880 2.800 ;
        RECT  3.475 0.490 3.710 0.925 ;
        RECT  2.025 0.695 3.475 0.925 ;
        RECT  3.190 1.155 3.390 1.385 ;
        RECT  2.960 1.155 3.190 2.800 ;
        RECT  2.285 2.565 2.515 3.375 ;
        RECT  2.025 2.565 2.285 2.795 ;
        RECT  1.795 0.470 2.025 2.795 ;
        RECT  1.255 0.975 1.485 2.655 ;
        RECT  0.180 0.975 1.255 1.205 ;
        RECT  0.180 2.425 1.255 2.655 ;
    END
END DFKSND2BWP7T

MACRO DFNCND0BWP7T
    CLASS CORE ;
    FOREIGN DFNCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.340 1.195 11.620 2.560 ;
        RECT  11.205 1.195 11.340 1.425 ;
        RECT  10.970 2.330 11.340 2.560 ;
        RECT  10.975 0.605 11.205 1.425 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.410 0.605 12.740 2.715 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4086 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.715 3.355 2.150 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 1.720 1.540 2.150 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.455 3.225 8.345 3.455 ;
        RECT  7.225 2.730 7.455 3.455 ;
        RECT  6.290 2.730 7.225 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.980 -0.235 12.880 0.235 ;
        RECT  11.640 -0.235 11.980 0.905 ;
        RECT  8.685 -0.235 11.640 0.235 ;
        RECT  8.345 -0.235 8.685 0.465 ;
        RECT  5.570 -0.235 8.345 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  0.520 -0.235 5.230 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.915 3.685 12.880 4.155 ;
        RECT  11.575 3.455 11.915 4.155 ;
        RECT  10.810 3.685 11.575 4.155 ;
        RECT  10.470 3.455 10.810 4.155 ;
        RECT  9.280 3.685 10.470 4.155 ;
        RECT  8.940 3.190 9.280 4.155 ;
        RECT  6.995 3.685 8.940 4.155 ;
        RECT  6.655 3.190 6.995 4.155 ;
        RECT  2.385 3.685 6.655 4.155 ;
        RECT  2.045 3.435 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.935 1.600 12.165 3.020 ;
        RECT  10.720 2.790 11.935 3.020 ;
        RECT  9.165 0.465 10.740 0.695 ;
        RECT  10.490 0.990 10.720 3.020 ;
        RECT  9.695 0.990 10.490 1.220 ;
        RECT  9.995 2.510 10.490 2.740 ;
        RECT  10.005 1.565 10.235 2.280 ;
        RECT  9.345 2.050 10.005 2.280 ;
        RECT  9.765 2.510 9.995 3.375 ;
        RECT  9.465 0.990 9.695 1.820 ;
        RECT  8.680 1.590 9.465 1.820 ;
        RECT  9.115 2.050 9.345 2.960 ;
        RECT  8.935 0.465 9.165 1.220 ;
        RECT  7.915 2.730 9.115 2.960 ;
        RECT  8.405 0.990 8.935 1.220 ;
        RECT  8.405 2.270 8.690 2.500 ;
        RECT  8.175 0.990 8.405 2.500 ;
        RECT  7.435 0.990 8.175 1.220 ;
        RECT  7.685 1.615 7.915 2.960 ;
        RECT  7.140 1.615 7.685 1.845 ;
        RECT  6.910 0.985 7.140 1.845 ;
        RECT  6.505 2.270 7.060 2.500 ;
        RECT  6.715 0.985 6.910 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.070 2.460 5.735 2.690 ;
        RECT  3.835 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  1.185 0.465 4.125 0.695 ;
        RECT  2.920 3.040 3.985 3.270 ;
        RECT  3.605 0.990 3.835 2.690 ;
        RECT  3.450 0.990 3.605 1.220 ;
        RECT  3.235 2.460 3.605 2.690 ;
        RECT  2.690 2.450 2.920 3.270 ;
        RECT  2.000 2.450 2.690 2.680 ;
        RECT  1.770 0.925 2.000 2.680 ;
        RECT  1.520 0.925 1.770 1.155 ;
        RECT  1.520 2.450 1.770 2.680 ;
        RECT  1.310 2.935 1.650 3.455 ;
        RECT  0.465 2.935 1.310 3.165 ;
        RECT  0.955 0.465 1.185 1.225 ;
        RECT  0.345 0.995 0.955 1.225 ;
        RECT  0.345 2.425 0.465 3.165 ;
        RECT  0.235 0.995 0.345 3.165 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFNCND0BWP7T

MACRO DFNCND1BWP7T
    CLASS CORE ;
    FOREIGN DFNCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.8520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.340 1.075 11.620 2.560 ;
        RECT  11.205 1.075 11.340 1.305 ;
        RECT  10.970 2.330 11.340 2.560 ;
        RECT  10.975 0.480 11.205 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.410 0.470 12.740 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4086 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.715 3.355 2.150 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 1.720 1.540 2.150 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.455 3.225 8.345 3.455 ;
        RECT  7.225 2.730 7.455 3.455 ;
        RECT  6.290 2.730 7.225 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.980 -0.235 12.880 0.235 ;
        RECT  11.640 -0.235 11.980 0.810 ;
        RECT  8.685 -0.235 11.640 0.235 ;
        RECT  8.345 -0.235 8.685 0.465 ;
        RECT  5.570 -0.235 8.345 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  0.520 -0.235 5.230 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.915 3.685 12.880 4.155 ;
        RECT  11.575 3.455 11.915 4.155 ;
        RECT  10.810 3.685 11.575 4.155 ;
        RECT  10.470 3.455 10.810 4.155 ;
        RECT  9.280 3.685 10.470 4.155 ;
        RECT  8.940 3.190 9.280 4.155 ;
        RECT  6.995 3.685 8.940 4.155 ;
        RECT  6.655 3.190 6.995 4.155 ;
        RECT  2.385 3.685 6.655 4.155 ;
        RECT  2.045 3.435 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.935 1.600 12.165 3.020 ;
        RECT  10.720 2.790 11.935 3.020 ;
        RECT  9.165 0.465 10.740 0.695 ;
        RECT  10.490 0.990 10.720 3.020 ;
        RECT  9.695 0.990 10.490 1.220 ;
        RECT  9.995 2.565 10.490 2.795 ;
        RECT  10.005 1.565 10.235 2.260 ;
        RECT  9.345 2.030 10.005 2.260 ;
        RECT  9.765 2.565 9.995 3.375 ;
        RECT  9.465 0.990 9.695 1.760 ;
        RECT  8.680 1.530 9.465 1.760 ;
        RECT  9.115 2.030 9.345 2.960 ;
        RECT  8.935 0.465 9.165 1.220 ;
        RECT  7.915 2.730 9.115 2.960 ;
        RECT  8.405 0.990 8.935 1.220 ;
        RECT  8.405 2.270 8.690 2.500 ;
        RECT  8.175 0.990 8.405 2.500 ;
        RECT  7.435 0.990 8.175 1.220 ;
        RECT  7.685 1.615 7.915 2.960 ;
        RECT  7.140 1.615 7.685 1.845 ;
        RECT  6.910 0.985 7.140 1.845 ;
        RECT  6.505 2.270 7.060 2.500 ;
        RECT  6.715 0.985 6.910 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.070 2.460 5.735 2.690 ;
        RECT  3.835 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  1.185 0.465 4.125 0.695 ;
        RECT  2.920 3.040 3.985 3.270 ;
        RECT  3.605 0.990 3.835 2.690 ;
        RECT  3.450 0.990 3.605 1.220 ;
        RECT  3.235 2.460 3.605 2.690 ;
        RECT  2.690 2.450 2.920 3.270 ;
        RECT  2.000 2.450 2.690 2.680 ;
        RECT  1.770 0.925 2.000 2.680 ;
        RECT  1.520 0.925 1.770 1.155 ;
        RECT  1.520 2.450 1.770 2.680 ;
        RECT  1.310 2.935 1.650 3.455 ;
        RECT  0.465 2.935 1.310 3.165 ;
        RECT  0.955 0.465 1.185 1.225 ;
        RECT  0.345 0.995 0.955 1.225 ;
        RECT  0.345 2.425 0.465 3.165 ;
        RECT  0.235 0.995 0.345 3.165 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFNCND1BWP7T

MACRO DFNCND2BWP7T
    CLASS CORE ;
    FOREIGN DFNCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.880 0.465 12.225 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.605 1.055 13.860 2.690 ;
        RECT  13.580 0.465 13.605 3.310 ;
        RECT  13.370 0.465 13.580 1.285 ;
        RECT  13.375 2.460 13.580 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4086 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.715 3.355 2.150 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.600 1.720 1.540 2.150 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.455 3.225 8.355 3.455 ;
        RECT  7.225 2.730 7.455 3.455 ;
        RECT  6.290 2.730 7.225 2.960 ;
        RECT  6.060 2.730 6.290 3.270 ;
        RECT  4.315 2.940 6.060 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 -0.235 14.560 0.235 ;
        RECT  14.095 -0.235 14.325 1.245 ;
        RECT  12.940 -0.235 14.095 0.235 ;
        RECT  12.600 -0.235 12.940 1.180 ;
        RECT  11.460 -0.235 12.600 0.235 ;
        RECT  11.120 -0.235 11.460 0.465 ;
        RECT  9.530 -0.235 11.120 0.235 ;
        RECT  9.190 -0.235 9.530 0.465 ;
        RECT  5.570 -0.235 9.190 0.235 ;
        RECT  5.230 -0.235 5.570 1.100 ;
        RECT  0.520 -0.235 5.230 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 3.685 14.560 4.155 ;
        RECT  14.095 2.255 14.325 4.155 ;
        RECT  12.940 3.685 14.095 4.155 ;
        RECT  12.600 3.250 12.940 4.155 ;
        RECT  11.345 3.685 12.600 4.155 ;
        RECT  11.005 3.250 11.345 4.155 ;
        RECT  9.745 3.685 11.005 4.155 ;
        RECT  9.405 3.190 9.745 4.155 ;
        RECT  6.995 3.685 9.405 4.155 ;
        RECT  6.655 3.190 6.995 4.155 ;
        RECT  2.385 3.685 6.655 4.155 ;
        RECT  2.045 3.435 2.385 4.155 ;
        RECT  1.080 3.685 2.045 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.895 1.600 13.125 3.020 ;
        RECT  11.120 2.790 12.895 3.020 ;
        RECT  11.410 0.695 11.640 1.940 ;
        RECT  8.715 0.695 11.410 0.925 ;
        RECT  10.890 1.155 11.120 3.020 ;
        RECT  9.675 1.155 10.890 1.385 ;
        RECT  10.465 2.540 10.890 2.770 ;
        RECT  10.360 1.670 10.590 2.260 ;
        RECT  10.235 2.540 10.465 3.370 ;
        RECT  9.695 2.030 10.360 2.260 ;
        RECT  9.465 2.030 9.695 2.960 ;
        RECT  9.445 1.155 9.675 1.750 ;
        RECT  7.915 2.730 9.465 2.960 ;
        RECT  8.945 1.520 9.445 1.750 ;
        RECT  8.715 2.270 8.910 2.500 ;
        RECT  8.485 0.465 8.715 2.500 ;
        RECT  7.435 0.990 8.485 1.220 ;
        RECT  7.685 1.615 7.915 2.960 ;
        RECT  7.140 1.615 7.685 1.845 ;
        RECT  6.910 0.985 7.140 1.845 ;
        RECT  6.505 2.270 7.060 2.500 ;
        RECT  6.715 0.985 6.910 1.220 ;
        RECT  6.280 1.330 6.505 2.500 ;
        RECT  6.275 0.870 6.280 2.500 ;
        RECT  6.050 0.870 6.275 1.560 ;
        RECT  5.250 1.330 6.050 1.560 ;
        RECT  5.585 1.790 5.925 2.230 ;
        RECT  4.070 2.460 5.735 2.690 ;
        RECT  3.835 2.000 5.585 2.230 ;
        RECT  4.910 1.330 5.250 1.770 ;
        RECT  1.185 0.465 4.125 0.695 ;
        RECT  2.920 3.040 3.985 3.270 ;
        RECT  3.605 0.990 3.835 2.690 ;
        RECT  3.450 0.990 3.605 1.220 ;
        RECT  3.235 2.460 3.605 2.690 ;
        RECT  2.690 2.450 2.920 3.270 ;
        RECT  2.000 2.450 2.690 2.680 ;
        RECT  1.770 0.925 2.000 2.680 ;
        RECT  1.520 0.925 1.770 1.155 ;
        RECT  1.520 2.450 1.770 2.680 ;
        RECT  1.310 2.935 1.650 3.455 ;
        RECT  0.465 2.935 1.310 3.165 ;
        RECT  0.955 0.465 1.185 1.225 ;
        RECT  0.345 0.995 0.955 1.225 ;
        RECT  0.345 2.425 0.465 3.165 ;
        RECT  0.235 0.995 0.345 3.165 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFNCND2BWP7T

MACRO DFND0BWP7T
    CLASS CORE ;
    FOREIGN DFND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.075 9.940 2.560 ;
        RECT  9.525 1.075 9.660 1.305 ;
        RECT  9.240 2.330 9.660 2.560 ;
        RECT  9.295 0.510 9.525 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.730 0.515 11.060 2.720 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.320 1.605 3.535 1.950 ;
        RECT  3.090 1.210 3.320 1.950 ;
        RECT  2.380 1.210 3.090 1.590 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 -0.235 11.200 0.235 ;
        RECT  9.960 -0.235 10.300 0.810 ;
        RECT  7.165 -0.235 9.960 0.235 ;
        RECT  6.825 -0.235 7.165 0.465 ;
        RECT  5.145 -0.235 6.825 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  0.520 -0.235 4.805 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.240 3.685 11.200 4.155 ;
        RECT  9.900 3.315 10.240 4.155 ;
        RECT  8.160 3.685 9.900 4.155 ;
        RECT  7.820 3.250 8.160 4.155 ;
        RECT  5.160 3.685 7.820 4.155 ;
        RECT  4.820 3.190 5.160 4.155 ;
        RECT  2.590 3.685 4.820 4.155 ;
        RECT  2.360 2.685 2.590 4.155 ;
        RECT  1.080 3.685 2.360 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.255 1.600 10.485 3.020 ;
        RECT  9.005 2.790 10.255 3.020 ;
        RECT  7.625 0.465 9.055 0.695 ;
        RECT  8.825 1.020 9.005 3.020 ;
        RECT  8.775 1.020 8.825 3.380 ;
        RECT  8.085 1.020 8.775 1.250 ;
        RECT  8.595 2.790 8.775 3.380 ;
        RECT  8.315 1.565 8.545 2.310 ;
        RECT  8.085 2.080 8.315 2.310 ;
        RECT  7.855 1.020 8.085 1.830 ;
        RECT  7.855 2.080 8.085 2.995 ;
        RECT  7.370 1.600 7.855 1.830 ;
        RECT  6.585 2.765 7.855 2.995 ;
        RECT  7.395 0.465 7.625 1.220 ;
        RECT  7.135 2.300 7.420 2.530 ;
        RECT  7.135 0.990 7.395 1.220 ;
        RECT  6.905 0.990 7.135 2.530 ;
        RECT  5.860 3.225 7.130 3.455 ;
        RECT  6.340 0.910 6.585 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.580 2.270 5.855 2.500 ;
        RECT  4.485 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.440 ;
        RECT  4.185 2.210 5.075 2.440 ;
        RECT  4.580 0.960 4.810 1.915 ;
        RECT  4.255 2.730 4.485 3.395 ;
        RECT  3.255 3.165 4.255 3.395 ;
        RECT  1.385 0.465 4.190 0.695 ;
        RECT  3.955 0.990 4.185 2.440 ;
        RECT  3.550 0.990 3.955 1.220 ;
        RECT  3.915 2.210 3.955 2.440 ;
        RECT  3.685 2.210 3.915 2.895 ;
        RECT  3.025 2.220 3.255 3.395 ;
        RECT  2.830 2.220 3.025 2.450 ;
        RECT  2.600 1.825 2.830 2.450 ;
        RECT  2.075 0.925 2.145 2.165 ;
        RECT  1.915 0.925 2.075 3.455 ;
        RECT  1.615 0.925 1.915 1.155 ;
        RECT  1.845 1.990 1.915 3.455 ;
        RECT  1.540 2.570 1.845 2.800 ;
        RECT  1.730 3.225 1.845 3.455 ;
        RECT  1.385 1.360 1.475 2.165 ;
        RECT  1.245 0.465 1.385 2.165 ;
        RECT  1.155 0.465 1.245 1.565 ;
        RECT  0.345 0.995 1.155 1.225 ;
        RECT  0.345 2.505 0.465 2.845 ;
        RECT  0.115 0.995 0.345 2.845 ;
    END
END DFND0BWP7T

MACRO DFND1BWP7T
    CLASS CORE ;
    FOREIGN DFND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.075 9.940 2.560 ;
        RECT  9.525 1.075 9.660 1.305 ;
        RECT  9.240 2.330 9.660 2.560 ;
        RECT  9.295 0.480 9.525 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.730 0.470 11.060 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.320 1.605 3.535 1.950 ;
        RECT  3.090 1.210 3.320 1.950 ;
        RECT  2.380 1.210 3.090 1.590 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 -0.235 11.200 0.235 ;
        RECT  9.960 -0.235 10.300 0.810 ;
        RECT  7.165 -0.235 9.960 0.235 ;
        RECT  6.825 -0.235 7.165 0.465 ;
        RECT  5.145 -0.235 6.825 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  0.520 -0.235 4.805 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 3.685 11.200 4.155 ;
        RECT  9.960 3.250 10.300 4.155 ;
        RECT  8.160 3.685 9.960 4.155 ;
        RECT  7.820 3.250 8.160 4.155 ;
        RECT  5.160 3.685 7.820 4.155 ;
        RECT  4.820 3.190 5.160 4.155 ;
        RECT  2.590 3.685 4.820 4.155 ;
        RECT  2.360 2.685 2.590 4.155 ;
        RECT  1.080 3.685 2.360 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.255 1.600 10.485 3.020 ;
        RECT  9.005 2.790 10.255 3.020 ;
        RECT  7.625 0.465 9.055 0.695 ;
        RECT  8.825 1.020 9.005 3.020 ;
        RECT  8.775 1.020 8.825 3.380 ;
        RECT  8.085 1.020 8.775 1.250 ;
        RECT  8.595 2.565 8.775 3.380 ;
        RECT  8.315 1.565 8.545 2.310 ;
        RECT  8.085 2.080 8.315 2.310 ;
        RECT  7.855 1.020 8.085 1.830 ;
        RECT  7.855 2.080 8.085 2.995 ;
        RECT  7.370 1.600 7.855 1.830 ;
        RECT  6.585 2.765 7.855 2.995 ;
        RECT  7.395 0.465 7.625 1.220 ;
        RECT  7.135 2.300 7.420 2.530 ;
        RECT  7.135 0.990 7.395 1.220 ;
        RECT  6.905 0.990 7.135 2.530 ;
        RECT  5.860 3.225 7.130 3.455 ;
        RECT  6.340 0.910 6.585 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.580 2.270 5.855 2.500 ;
        RECT  4.485 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.440 ;
        RECT  4.185 2.210 5.075 2.440 ;
        RECT  4.580 0.960 4.810 1.915 ;
        RECT  4.255 2.730 4.485 3.395 ;
        RECT  3.255 3.165 4.255 3.395 ;
        RECT  1.385 0.465 4.190 0.695 ;
        RECT  3.955 0.990 4.185 2.440 ;
        RECT  3.550 0.990 3.955 1.220 ;
        RECT  3.915 2.210 3.955 2.440 ;
        RECT  3.685 2.210 3.915 2.895 ;
        RECT  3.025 2.220 3.255 3.395 ;
        RECT  2.830 2.220 3.025 2.450 ;
        RECT  2.600 1.825 2.830 2.450 ;
        RECT  2.075 0.925 2.145 2.165 ;
        RECT  1.915 0.925 2.075 3.455 ;
        RECT  1.615 0.925 1.915 1.155 ;
        RECT  1.845 1.990 1.915 3.455 ;
        RECT  1.540 2.570 1.845 2.800 ;
        RECT  1.730 3.225 1.845 3.455 ;
        RECT  1.385 1.360 1.475 2.165 ;
        RECT  1.245 0.465 1.385 2.165 ;
        RECT  1.155 0.465 1.245 1.565 ;
        RECT  0.345 0.995 1.155 1.225 ;
        RECT  0.345 2.505 0.465 2.845 ;
        RECT  0.115 0.995 0.345 2.845 ;
    END
END DFND1BWP7T

MACRO DFND2BWP7T
    CLASS CORE ;
    FOREIGN DFND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.200 0.465 10.545 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.925 1.055 12.180 2.690 ;
        RECT  11.900 0.465 11.925 3.310 ;
        RECT  11.690 0.465 11.900 1.285 ;
        RECT  11.695 2.460 11.900 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.320 1.605 3.535 1.950 ;
        RECT  3.090 1.210 3.320 1.950 ;
        RECT  2.380 1.210 3.090 1.590 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 -0.235 12.880 0.235 ;
        RECT  12.415 -0.235 12.645 1.245 ;
        RECT  11.260 -0.235 12.415 0.235 ;
        RECT  10.920 -0.235 11.260 1.180 ;
        RECT  9.780 -0.235 10.920 0.235 ;
        RECT  9.440 -0.235 9.780 0.465 ;
        RECT  8.165 -0.235 9.440 0.235 ;
        RECT  7.825 -0.235 8.165 0.465 ;
        RECT  5.145 -0.235 7.825 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  0.520 -0.235 4.805 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 3.685 12.880 4.155 ;
        RECT  12.415 2.255 12.645 4.155 ;
        RECT  11.260 3.685 12.415 4.155 ;
        RECT  10.920 3.250 11.260 4.155 ;
        RECT  9.780 3.685 10.920 4.155 ;
        RECT  9.440 3.250 9.780 4.155 ;
        RECT  8.165 3.685 9.440 4.155 ;
        RECT  7.825 3.250 8.165 4.155 ;
        RECT  5.160 3.685 7.825 4.155 ;
        RECT  4.820 3.190 5.160 4.155 ;
        RECT  2.590 3.685 4.820 4.155 ;
        RECT  2.360 2.685 2.590 4.155 ;
        RECT  1.080 3.685 2.360 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.215 1.605 11.445 3.010 ;
        RECT  9.365 2.780 11.215 3.010 ;
        RECT  9.730 0.695 9.960 1.945 ;
        RECT  7.645 0.695 9.730 0.925 ;
        RECT  9.135 1.155 9.365 3.010 ;
        RECT  8.235 1.155 9.135 1.385 ;
        RECT  8.940 2.565 9.135 3.010 ;
        RECT  8.710 2.565 8.940 3.380 ;
        RECT  8.600 1.675 8.830 2.310 ;
        RECT  8.185 2.080 8.600 2.310 ;
        RECT  8.005 1.155 8.235 1.830 ;
        RECT  7.955 2.080 8.185 2.995 ;
        RECT  7.380 1.600 8.005 1.830 ;
        RECT  6.585 2.765 7.955 2.995 ;
        RECT  7.415 0.695 7.645 1.220 ;
        RECT  7.115 2.300 7.420 2.530 ;
        RECT  7.115 0.990 7.415 1.220 ;
        RECT  6.885 0.990 7.115 2.530 ;
        RECT  5.860 3.225 7.020 3.455 ;
        RECT  6.340 0.910 6.585 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.580 2.270 5.855 2.500 ;
        RECT  4.485 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.440 ;
        RECT  4.185 2.210 5.075 2.440 ;
        RECT  4.580 0.960 4.810 1.915 ;
        RECT  4.255 2.730 4.485 3.395 ;
        RECT  3.255 3.165 4.255 3.395 ;
        RECT  1.385 0.465 4.190 0.695 ;
        RECT  3.955 0.990 4.185 2.440 ;
        RECT  3.550 0.990 3.955 1.220 ;
        RECT  3.915 2.210 3.955 2.440 ;
        RECT  3.685 2.210 3.915 2.895 ;
        RECT  3.025 2.220 3.255 3.395 ;
        RECT  2.830 2.220 3.025 2.450 ;
        RECT  2.600 1.825 2.830 2.450 ;
        RECT  2.075 0.925 2.145 2.165 ;
        RECT  1.915 0.925 2.075 3.455 ;
        RECT  1.615 0.925 1.915 1.155 ;
        RECT  1.845 1.990 1.915 3.455 ;
        RECT  1.540 2.570 1.845 2.800 ;
        RECT  1.730 3.225 1.845 3.455 ;
        RECT  1.385 1.360 1.475 2.165 ;
        RECT  1.245 0.465 1.385 2.165 ;
        RECT  1.155 0.465 1.245 1.565 ;
        RECT  0.345 0.995 1.155 1.225 ;
        RECT  0.345 2.505 0.465 2.845 ;
        RECT  0.115 0.995 0.345 2.845 ;
    END
END DFND2BWP7T

MACRO DFNSND0BWP7T
    CLASS CORE ;
    FOREIGN DFNSND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.970 0.515 13.300 2.715 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.075 12.180 2.665 ;
        RECT  11.765 1.075 11.900 1.305 ;
        RECT  11.480 2.435 11.900 2.665 ;
        RECT  11.535 0.510 11.765 1.305 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4086 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.700 3.460 2.150 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 -0.235 13.440 0.235 ;
        RECT  12.200 -0.235 12.540 0.810 ;
        RECT  10.210 -0.235 12.200 0.235 ;
        RECT  9.870 -0.235 10.210 0.950 ;
        RECT  5.170 -0.235 9.870 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  0.520 -0.235 4.830 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.460 3.685 13.440 4.155 ;
        RECT  12.120 3.455 12.460 4.155 ;
        RECT  10.355 3.685 12.120 4.155 ;
        RECT  10.015 3.455 10.355 4.155 ;
        RECT  9.330 3.685 10.015 4.155 ;
        RECT  8.990 3.450 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.995 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.495 1.600 12.725 3.225 ;
        RECT  10.230 2.995 12.495 3.225 ;
        RECT  11.250 1.635 11.670 1.865 ;
        RECT  11.065 0.720 11.250 2.230 ;
        RECT  11.020 0.720 11.065 2.690 ;
        RECT  10.630 0.720 11.020 0.950 ;
        RECT  10.835 2.000 11.020 2.690 ;
        RECT  9.720 2.000 10.835 2.230 ;
        RECT  10.385 1.205 10.730 1.770 ;
        RECT  9.440 1.205 10.385 1.435 ;
        RECT  9.995 2.465 10.230 3.225 ;
        RECT  8.485 2.465 9.995 2.695 ;
        RECT  9.380 1.780 9.720 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.630 ;
        RECT  1.130 0.465 4.130 0.695 ;
        RECT  3.150 3.040 4.120 3.270 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.400 3.920 2.630 ;
        RECT  2.920 2.525 3.150 3.270 ;
        RECT  2.045 2.525 2.920 2.755 ;
        RECT  1.815 0.925 2.045 2.755 ;
        RECT  1.520 0.925 1.815 1.155 ;
        RECT  1.520 2.525 1.815 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.900 0.465 1.130 1.210 ;
        RECT  0.345 0.980 0.900 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFNSND0BWP7T

MACRO DFNSND1BWP7T
    CLASS CORE ;
    FOREIGN DFNSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.970 0.470 13.300 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.075 12.180 2.560 ;
        RECT  11.765 1.075 11.900 1.305 ;
        RECT  11.480 2.330 11.900 2.560 ;
        RECT  11.535 0.465 11.765 1.305 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4086 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.700 3.460 2.150 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 -0.235 13.440 0.235 ;
        RECT  12.200 -0.235 12.540 0.810 ;
        RECT  10.210 -0.235 12.200 0.235 ;
        RECT  9.870 -0.235 10.210 0.930 ;
        RECT  5.170 -0.235 9.870 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  0.520 -0.235 4.830 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 3.685 13.440 4.155 ;
        RECT  12.200 3.250 12.540 4.155 ;
        RECT  10.355 3.685 12.200 4.155 ;
        RECT  10.015 3.455 10.355 4.155 ;
        RECT  9.330 3.685 10.015 4.155 ;
        RECT  8.990 3.450 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.995 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.495 1.600 12.725 3.020 ;
        RECT  11.725 2.790 12.495 3.020 ;
        RECT  11.495 2.790 11.725 3.225 ;
        RECT  11.250 1.635 11.670 1.865 ;
        RECT  10.230 2.995 11.495 3.225 ;
        RECT  11.065 0.680 11.250 2.230 ;
        RECT  11.020 0.680 11.065 2.765 ;
        RECT  10.630 0.680 11.020 0.910 ;
        RECT  10.835 2.000 11.020 2.765 ;
        RECT  9.720 2.000 10.835 2.230 ;
        RECT  10.385 1.205 10.730 1.770 ;
        RECT  9.440 1.205 10.385 1.435 ;
        RECT  9.995 2.465 10.230 3.225 ;
        RECT  8.485 2.465 9.995 2.695 ;
        RECT  9.380 1.780 9.720 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.630 ;
        RECT  1.130 0.465 4.130 0.695 ;
        RECT  3.150 3.040 4.120 3.270 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.400 3.920 2.630 ;
        RECT  2.920 2.525 3.150 3.270 ;
        RECT  2.045 2.525 2.920 2.755 ;
        RECT  1.815 0.925 2.045 2.755 ;
        RECT  1.520 0.925 1.815 1.155 ;
        RECT  1.520 2.525 1.815 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.900 0.465 1.130 1.210 ;
        RECT  0.345 0.980 0.900 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFNSND1BWP7T

MACRO DFNSND2BWP7T
    CLASS CORE ;
    FOREIGN DFNSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.165 1.055 14.420 2.730 ;
        RECT  14.140 0.470 14.165 3.310 ;
        RECT  13.935 0.470 14.140 1.290 ;
        RECT  13.935 2.500 14.140 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.440 0.510 12.780 2.560 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4086 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.700 3.460 2.150 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.885 -0.235 15.120 0.235 ;
        RECT  14.655 -0.235 14.885 1.290 ;
        RECT  13.500 -0.235 14.655 0.235 ;
        RECT  13.160 -0.235 13.500 1.205 ;
        RECT  11.995 -0.235 13.160 0.235 ;
        RECT  11.655 -0.235 11.995 1.205 ;
        RECT  10.345 -0.235 11.655 0.235 ;
        RECT  10.005 -0.235 10.345 0.930 ;
        RECT  5.170 -0.235 10.005 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  0.520 -0.235 4.830 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.885 3.685 15.120 4.155 ;
        RECT  14.655 2.255 14.885 4.155 ;
        RECT  13.500 3.685 14.655 4.155 ;
        RECT  13.160 3.250 13.500 4.155 ;
        RECT  11.930 3.685 13.160 4.155 ;
        RECT  11.590 3.455 11.930 4.155 ;
        RECT  10.450 3.685 11.590 4.155 ;
        RECT  10.110 3.455 10.450 4.155 ;
        RECT  9.330 3.685 10.110 4.155 ;
        RECT  8.990 3.225 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.995 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.455 1.600 13.685 3.020 ;
        RECT  12.285 2.790 13.455 3.020 ;
        RECT  12.055 2.790 12.285 3.225 ;
        RECT  11.370 1.635 12.210 1.865 ;
        RECT  10.245 2.995 12.055 3.225 ;
        RECT  11.160 0.680 11.370 2.230 ;
        RECT  11.140 0.680 11.160 2.765 ;
        RECT  10.765 0.680 11.140 0.910 ;
        RECT  10.930 2.000 11.140 2.765 ;
        RECT  9.815 2.000 10.930 2.230 ;
        RECT  10.480 1.205 10.865 1.770 ;
        RECT  9.440 1.205 10.480 1.435 ;
        RECT  10.010 2.465 10.245 3.225 ;
        RECT  8.485 2.465 10.010 2.695 ;
        RECT  9.475 1.780 9.815 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.630 ;
        RECT  1.130 0.465 4.130 0.695 ;
        RECT  3.150 3.040 4.120 3.270 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.400 3.920 2.630 ;
        RECT  2.920 2.525 3.150 3.270 ;
        RECT  2.045 2.525 2.920 2.755 ;
        RECT  1.815 0.925 2.045 2.755 ;
        RECT  1.520 0.925 1.815 1.155 ;
        RECT  1.520 2.525 1.815 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.900 0.465 1.130 1.210 ;
        RECT  0.345 0.980 0.900 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFNSND2BWP7T

MACRO DFQD0BWP7T
    CLASS CORE ;
    FOREIGN DFQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.170 0.530 10.500 3.180 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 1.715 3.460 2.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 -0.235 10.640 0.235 ;
        RECT  9.430 -0.235 9.660 0.820 ;
        RECT  8.195 -0.235 9.430 0.235 ;
        RECT  7.855 -0.235 8.195 0.795 ;
        RECT  5.145 -0.235 7.855 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  2.560 -0.235 4.805 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.685 3.685 10.640 4.155 ;
        RECT  9.455 2.845 9.685 4.155 ;
        RECT  8.185 3.685 9.455 4.155 ;
        RECT  7.845 3.250 8.185 4.155 ;
        RECT  5.155 3.685 7.845 4.155 ;
        RECT  4.795 3.190 5.155 4.155 ;
        RECT  2.590 3.685 4.795 4.155 ;
        RECT  2.250 2.800 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.185 1.650 9.930 1.890 ;
        RECT  8.955 1.065 9.185 3.340 ;
        RECT  8.865 1.065 8.955 1.295 ;
        RECT  8.620 3.110 8.955 3.340 ;
        RECT  8.635 0.510 8.865 1.295 ;
        RECT  8.415 1.565 8.645 2.340 ;
        RECT  8.085 1.065 8.635 1.295 ;
        RECT  8.135 2.110 8.415 2.340 ;
        RECT  7.905 2.110 8.135 2.995 ;
        RECT  7.855 1.065 8.085 1.880 ;
        RECT  6.570 2.765 7.905 2.995 ;
        RECT  7.370 1.650 7.855 1.880 ;
        RECT  7.135 2.300 7.405 2.530 ;
        RECT  7.135 0.990 7.350 1.220 ;
        RECT  6.905 0.990 7.135 2.530 ;
        RECT  5.860 3.225 7.115 3.455 ;
        RECT  6.340 0.910 6.570 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.565 2.270 5.855 2.500 ;
        RECT  4.540 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.415 ;
        RECT  4.050 2.185 5.075 2.415 ;
        RECT  4.580 0.960 4.810 1.890 ;
        RECT  4.310 2.730 4.540 3.280 ;
        RECT  3.140 3.050 4.310 3.280 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.820 0.990 4.050 2.695 ;
        RECT  3.520 0.990 3.820 1.220 ;
        RECT  3.485 2.465 3.820 2.695 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.910 2.340 3.140 3.280 ;
        RECT  2.020 0.975 2.930 1.205 ;
        RECT  2.020 2.340 2.910 2.570 ;
        RECT  1.790 0.975 2.020 2.755 ;
        RECT  1.520 0.975 1.790 1.205 ;
        RECT  1.520 2.525 1.790 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.995 0.530 1.225 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.995 0.345 3.215 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFQD0BWP7T

MACRO DFQD1BWP7T
    CLASS CORE ;
    FOREIGN DFQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.170 0.470 10.500 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 1.715 3.460 2.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 -0.235 10.640 0.235 ;
        RECT  9.430 -0.235 9.660 1.270 ;
        RECT  8.195 -0.235 9.430 0.235 ;
        RECT  7.855 -0.235 8.195 0.770 ;
        RECT  5.145 -0.235 7.855 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  2.560 -0.235 4.805 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.685 3.685 10.640 4.155 ;
        RECT  9.455 2.255 9.685 4.155 ;
        RECT  8.185 3.685 9.455 4.155 ;
        RECT  7.845 3.250 8.185 4.155 ;
        RECT  5.155 3.685 7.845 4.155 ;
        RECT  4.795 3.190 5.155 4.155 ;
        RECT  2.590 3.685 4.795 4.155 ;
        RECT  2.250 2.800 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.185 1.650 9.930 1.890 ;
        RECT  8.955 1.020 9.185 2.805 ;
        RECT  8.865 1.020 8.955 1.250 ;
        RECT  8.905 2.565 8.955 2.805 ;
        RECT  8.675 2.565 8.905 3.380 ;
        RECT  8.635 0.495 8.865 1.250 ;
        RECT  8.085 1.020 8.635 1.250 ;
        RECT  8.395 1.565 8.625 2.340 ;
        RECT  8.135 2.110 8.395 2.340 ;
        RECT  7.905 2.110 8.135 2.995 ;
        RECT  7.855 1.020 8.085 1.880 ;
        RECT  6.570 2.765 7.905 2.995 ;
        RECT  7.370 1.650 7.855 1.880 ;
        RECT  7.135 2.300 7.405 2.530 ;
        RECT  7.135 0.990 7.350 1.220 ;
        RECT  6.905 0.990 7.135 2.530 ;
        RECT  5.860 3.225 7.115 3.455 ;
        RECT  6.340 0.910 6.570 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.565 2.270 5.855 2.500 ;
        RECT  4.540 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.415 ;
        RECT  4.050 2.185 5.075 2.415 ;
        RECT  4.580 0.960 4.810 1.890 ;
        RECT  4.310 2.730 4.540 3.280 ;
        RECT  3.140 3.050 4.310 3.280 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.820 0.990 4.050 2.695 ;
        RECT  3.520 0.990 3.820 1.220 ;
        RECT  3.485 2.465 3.820 2.695 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.910 2.340 3.140 3.280 ;
        RECT  2.020 0.975 2.930 1.205 ;
        RECT  2.020 2.340 2.910 2.570 ;
        RECT  1.790 0.975 2.020 2.755 ;
        RECT  1.520 0.975 1.790 1.205 ;
        RECT  1.520 2.525 1.790 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.995 0.530 1.225 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.995 0.345 3.215 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFQD1BWP7T

MACRO DFQD2BWP7T
    CLASS CORE ;
    FOREIGN DFQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.245 1.055 10.500 2.730 ;
        RECT  10.220 0.470 10.245 3.310 ;
        RECT  10.015 0.470 10.220 1.290 ;
        RECT  10.015 2.500 10.220 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 1.715 3.460 2.110 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.965 -0.235 11.200 0.235 ;
        RECT  10.735 -0.235 10.965 1.270 ;
        RECT  9.500 -0.235 10.735 0.235 ;
        RECT  9.270 -0.235 9.500 1.270 ;
        RECT  8.130 -0.235 9.270 0.235 ;
        RECT  7.790 -0.235 8.130 0.770 ;
        RECT  5.145 -0.235 7.790 0.235 ;
        RECT  4.805 -0.235 5.145 0.730 ;
        RECT  2.560 -0.235 4.805 0.235 ;
        RECT  2.220 -0.235 2.560 0.730 ;
        RECT  0.520 -0.235 2.220 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.965 3.685 11.200 4.155 ;
        RECT  10.735 2.255 10.965 4.155 ;
        RECT  9.525 3.685 10.735 4.155 ;
        RECT  9.295 2.255 9.525 4.155 ;
        RECT  8.160 3.685 9.295 4.155 ;
        RECT  7.820 3.250 8.160 4.155 ;
        RECT  5.155 3.685 7.820 4.155 ;
        RECT  4.795 3.190 5.155 4.155 ;
        RECT  2.590 3.685 4.795 4.155 ;
        RECT  2.250 2.800 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.040 1.650 9.985 1.890 ;
        RECT  8.825 1.020 9.040 2.825 ;
        RECT  8.810 1.020 8.825 3.400 ;
        RECT  8.800 1.020 8.810 1.250 ;
        RECT  8.595 2.585 8.810 3.400 ;
        RECT  8.570 0.495 8.800 1.250 ;
        RECT  7.955 1.020 8.570 1.250 ;
        RECT  8.330 1.565 8.560 2.340 ;
        RECT  8.135 2.110 8.330 2.340 ;
        RECT  7.905 2.110 8.135 2.995 ;
        RECT  7.725 1.020 7.955 1.880 ;
        RECT  6.570 2.765 7.905 2.995 ;
        RECT  7.370 1.650 7.725 1.880 ;
        RECT  7.135 2.300 7.405 2.530 ;
        RECT  7.135 0.990 7.350 1.220 ;
        RECT  6.905 0.990 7.135 2.530 ;
        RECT  5.860 3.225 7.115 3.455 ;
        RECT  6.340 0.910 6.570 2.995 ;
        RECT  5.855 0.960 6.085 2.500 ;
        RECT  5.630 2.730 5.860 3.455 ;
        RECT  4.810 0.960 5.855 1.190 ;
        RECT  5.565 2.270 5.855 2.500 ;
        RECT  4.540 2.730 5.630 2.960 ;
        RECT  5.305 1.560 5.610 1.900 ;
        RECT  5.075 1.560 5.305 2.415 ;
        RECT  4.050 2.185 5.075 2.415 ;
        RECT  4.580 0.960 4.810 1.890 ;
        RECT  4.310 2.730 4.540 3.280 ;
        RECT  3.140 3.050 4.310 3.280 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.820 0.990 4.050 2.695 ;
        RECT  3.520 0.990 3.820 1.220 ;
        RECT  3.485 2.465 3.820 2.695 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.910 2.340 3.140 3.280 ;
        RECT  2.020 0.975 2.930 1.205 ;
        RECT  2.020 2.340 2.910 2.570 ;
        RECT  1.790 0.975 2.020 2.755 ;
        RECT  1.520 0.975 1.790 1.205 ;
        RECT  1.520 2.525 1.790 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.995 0.530 1.225 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.995 0.345 3.215 ;
        RECT  0.115 0.995 0.235 2.765 ;
    END
END DFQD2BWP7T

MACRO DFSND0BWP7T
    CLASS CORE ;
    FOREIGN DFSND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.970 0.515 13.300 2.715 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.075 12.180 2.665 ;
        RECT  11.765 1.075 11.900 1.305 ;
        RECT  11.480 2.435 11.900 2.665 ;
        RECT  11.535 0.510 11.765 1.305 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.715 3.460 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 -0.235 13.440 0.235 ;
        RECT  12.200 -0.235 12.540 0.810 ;
        RECT  10.210 -0.235 12.200 0.235 ;
        RECT  9.870 -0.235 10.210 0.950 ;
        RECT  5.170 -0.235 9.870 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  2.580 -0.235 4.830 0.235 ;
        RECT  2.240 -0.235 2.580 0.730 ;
        RECT  0.520 -0.235 2.240 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.460 3.685 13.440 4.155 ;
        RECT  12.120 3.455 12.460 4.155 ;
        RECT  10.355 3.685 12.120 4.155 ;
        RECT  10.015 3.455 10.355 4.155 ;
        RECT  9.330 3.685 10.015 4.155 ;
        RECT  8.990 3.455 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.330 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.495 1.540 12.725 3.225 ;
        RECT  10.230 2.995 12.495 3.225 ;
        RECT  11.250 1.635 11.670 1.865 ;
        RECT  11.065 0.720 11.250 2.230 ;
        RECT  11.020 0.720 11.065 2.690 ;
        RECT  10.630 0.720 11.020 0.950 ;
        RECT  10.835 2.000 11.020 2.690 ;
        RECT  9.720 2.000 10.835 2.230 ;
        RECT  10.385 1.205 10.730 1.770 ;
        RECT  9.440 1.205 10.385 1.435 ;
        RECT  9.995 2.465 10.230 3.225 ;
        RECT  8.485 2.465 9.995 2.695 ;
        RECT  9.380 1.780 9.720 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.640 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.410 3.920 2.640 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.005 0.975 2.930 1.205 ;
        RECT  1.775 0.975 2.005 2.755 ;
        RECT  1.520 0.975 1.775 1.205 ;
        RECT  1.520 2.525 1.775 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.980 0.530 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFSND0BWP7T

MACRO DFSND1BWP7T
    CLASS CORE ;
    FOREIGN DFSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.970 0.470 13.300 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.075 12.180 2.560 ;
        RECT  11.765 1.075 11.900 1.305 ;
        RECT  11.480 2.330 11.900 2.560 ;
        RECT  11.535 0.465 11.765 1.305 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.715 3.460 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 -0.235 13.440 0.235 ;
        RECT  12.200 -0.235 12.540 0.810 ;
        RECT  10.210 -0.235 12.200 0.235 ;
        RECT  9.870 -0.235 10.210 0.930 ;
        RECT  5.170 -0.235 9.870 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  2.580 -0.235 4.830 0.235 ;
        RECT  2.240 -0.235 2.580 0.730 ;
        RECT  0.520 -0.235 2.240 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 3.685 13.440 4.155 ;
        RECT  12.200 3.250 12.540 4.155 ;
        RECT  10.355 3.685 12.200 4.155 ;
        RECT  10.015 3.455 10.355 4.155 ;
        RECT  9.330 3.685 10.015 4.155 ;
        RECT  8.990 3.450 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.330 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.495 1.600 12.725 3.020 ;
        RECT  11.725 2.790 12.495 3.020 ;
        RECT  11.495 2.790 11.725 3.225 ;
        RECT  11.250 1.635 11.670 1.865 ;
        RECT  9.965 2.995 11.495 3.225 ;
        RECT  11.065 0.680 11.250 2.230 ;
        RECT  11.020 0.680 11.065 2.765 ;
        RECT  10.630 0.680 11.020 0.910 ;
        RECT  10.835 2.000 11.020 2.765 ;
        RECT  9.720 2.000 10.835 2.230 ;
        RECT  10.385 1.205 10.730 1.770 ;
        RECT  9.440 1.205 10.385 1.435 ;
        RECT  9.730 2.465 9.965 3.225 ;
        RECT  8.485 2.465 9.730 2.695 ;
        RECT  9.380 1.780 9.720 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.640 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.410 3.920 2.640 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.005 0.975 2.930 1.205 ;
        RECT  1.775 0.975 2.005 2.755 ;
        RECT  1.520 0.975 1.775 1.205 ;
        RECT  1.520 2.525 1.775 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.980 0.530 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFSND1BWP7T

MACRO DFSND2BWP7T
    CLASS CORE ;
    FOREIGN DFSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.165 1.055 14.420 2.730 ;
        RECT  14.140 0.470 14.165 3.310 ;
        RECT  13.935 0.470 14.140 1.290 ;
        RECT  13.935 2.500 14.140 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.440 0.510 12.780 2.560 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.715 3.460 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.885 -0.235 15.120 0.235 ;
        RECT  14.655 -0.235 14.885 1.290 ;
        RECT  13.500 -0.235 14.655 0.235 ;
        RECT  13.160 -0.235 13.500 1.205 ;
        RECT  11.995 -0.235 13.160 0.235 ;
        RECT  11.655 -0.235 11.995 1.205 ;
        RECT  10.345 -0.235 11.655 0.235 ;
        RECT  10.005 -0.235 10.345 0.930 ;
        RECT  5.170 -0.235 10.005 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  2.580 -0.235 4.830 0.235 ;
        RECT  2.240 -0.235 2.580 0.730 ;
        RECT  0.520 -0.235 2.240 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.885 3.685 15.120 4.155 ;
        RECT  14.655 2.255 14.885 4.155 ;
        RECT  13.500 3.685 14.655 4.155 ;
        RECT  13.160 3.250 13.500 4.155 ;
        RECT  11.930 3.685 13.160 4.155 ;
        RECT  11.590 3.455 11.930 4.155 ;
        RECT  10.450 3.685 11.590 4.155 ;
        RECT  10.110 3.455 10.450 4.155 ;
        RECT  9.330 3.685 10.110 4.155 ;
        RECT  8.990 3.225 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.330 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.455 1.600 13.685 3.020 ;
        RECT  12.285 2.790 13.455 3.020 ;
        RECT  12.055 2.790 12.285 3.225 ;
        RECT  11.370 1.635 12.210 1.865 ;
        RECT  10.245 2.995 12.055 3.225 ;
        RECT  11.160 0.680 11.370 2.230 ;
        RECT  11.140 0.680 11.160 2.765 ;
        RECT  10.765 0.680 11.140 0.910 ;
        RECT  10.930 2.000 11.140 2.765 ;
        RECT  9.815 2.000 10.930 2.230 ;
        RECT  10.480 1.205 10.865 1.770 ;
        RECT  9.440 1.205 10.480 1.435 ;
        RECT  10.010 2.465 10.245 3.225 ;
        RECT  8.485 2.465 10.010 2.695 ;
        RECT  9.475 1.780 9.815 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.640 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.410 3.920 2.640 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.005 0.975 2.930 1.205 ;
        RECT  1.775 0.975 2.005 2.755 ;
        RECT  1.520 0.975 1.775 1.205 ;
        RECT  1.520 2.525 1.775 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.980 0.530 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFSND2BWP7T

MACRO DFSNQD1BWP7T
    CLASS CORE ;
    FOREIGN DFSNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.925 1.075 12.180 2.560 ;
        RECT  11.900 0.465 11.925 3.265 ;
        RECT  11.695 0.465 11.900 1.305 ;
        RECT  11.695 2.330 11.900 3.265 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.715 3.460 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 -0.235 12.880 0.235 ;
        RECT  12.415 -0.235 12.645 1.240 ;
        RECT  10.210 -0.235 12.415 0.235 ;
        RECT  9.870 -0.235 10.210 0.930 ;
        RECT  5.170 -0.235 9.870 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  2.580 -0.235 4.830 0.235 ;
        RECT  2.240 -0.235 2.580 0.730 ;
        RECT  0.520 -0.235 2.240 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.645 3.685 12.880 4.155 ;
        RECT  12.415 2.255 12.645 4.155 ;
        RECT  10.560 3.685 12.415 4.155 ;
        RECT  10.220 2.545 10.560 4.155 ;
        RECT  9.330 3.685 10.220 4.155 ;
        RECT  8.990 3.260 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.330 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.225 1.635 11.670 1.865 ;
        RECT  10.995 0.680 11.225 3.305 ;
        RECT  10.690 0.680 10.995 0.910 ;
        RECT  9.720 2.000 10.995 2.230 ;
        RECT  10.385 1.205 10.730 1.770 ;
        RECT  9.440 1.205 10.385 1.435 ;
        RECT  8.485 2.465 9.815 2.695 ;
        RECT  9.380 1.780 9.720 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.640 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.410 3.920 2.640 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.005 0.975 2.930 1.205 ;
        RECT  1.775 0.975 2.005 2.755 ;
        RECT  1.520 0.975 1.775 1.205 ;
        RECT  1.520 2.525 1.775 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.980 0.530 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFSNQD1BWP7T

MACRO DFSNQD2BWP7T
    CLASS CORE ;
    FOREIGN DFSNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.940 8.695 3.340 ;
        RECT  7.125 2.940 8.355 3.220 ;
        RECT  6.895 2.730 7.125 3.220 ;
        RECT  5.370 2.730 6.895 2.960 ;
        RECT  5.140 2.730 5.370 3.155 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.485 1.040 12.740 2.740 ;
        RECT  12.460 0.465 12.485 3.325 ;
        RECT  12.255 0.465 12.460 1.275 ;
        RECT  12.255 2.510 12.460 3.325 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3348 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.715 3.460 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.700 1.540 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.205 -0.235 13.440 0.235 ;
        RECT  12.975 -0.235 13.205 1.240 ;
        RECT  11.765 -0.235 12.975 0.235 ;
        RECT  11.535 -0.235 11.765 1.240 ;
        RECT  10.210 -0.235 11.535 0.235 ;
        RECT  9.870 -0.235 10.210 0.930 ;
        RECT  5.170 -0.235 9.870 0.235 ;
        RECT  4.830 -0.235 5.170 0.960 ;
        RECT  2.580 -0.235 4.830 0.235 ;
        RECT  2.240 -0.235 2.580 0.730 ;
        RECT  0.520 -0.235 2.240 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.205 3.685 13.440 4.155 ;
        RECT  12.975 2.255 13.205 4.155 ;
        RECT  11.765 3.685 12.975 4.155 ;
        RECT  11.535 2.255 11.765 4.155 ;
        RECT  10.350 3.685 11.535 4.155 ;
        RECT  10.010 3.455 10.350 4.155 ;
        RECT  9.330 3.685 10.010 4.155 ;
        RECT  8.990 3.260 9.330 4.155 ;
        RECT  6.560 3.685 8.990 4.155 ;
        RECT  6.220 3.190 6.560 4.155 ;
        RECT  4.850 3.685 6.220 4.155 ;
        RECT  4.620 3.130 4.850 4.155 ;
        RECT  2.590 3.685 4.620 4.155 ;
        RECT  2.250 2.330 2.590 4.155 ;
        RECT  1.080 3.685 2.250 4.155 ;
        RECT  0.740 3.455 1.080 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.225 1.660 12.230 1.890 ;
        RECT  11.065 0.680 11.225 2.230 ;
        RECT  10.995 0.680 11.065 3.305 ;
        RECT  10.705 0.680 10.995 0.910 ;
        RECT  10.835 2.000 10.995 3.305 ;
        RECT  9.720 2.000 10.835 2.230 ;
        RECT  10.385 1.205 10.730 1.770 ;
        RECT  9.440 1.205 10.385 1.435 ;
        RECT  8.485 2.465 9.815 2.695 ;
        RECT  9.380 1.780 9.720 2.230 ;
        RECT  9.210 0.465 9.440 1.435 ;
        RECT  7.220 0.465 9.210 0.695 ;
        RECT  8.485 0.990 8.810 1.220 ;
        RECT  8.255 0.990 8.485 2.695 ;
        RECT  7.655 0.990 8.255 1.220 ;
        RECT  7.535 1.615 7.765 2.585 ;
        RECT  7.220 1.615 7.535 1.845 ;
        RECT  6.990 0.465 7.220 1.845 ;
        RECT  6.670 2.270 7.100 2.500 ;
        RECT  6.440 0.935 6.670 2.500 ;
        RECT  6.150 0.935 6.440 1.165 ;
        RECT  4.835 2.270 6.440 2.500 ;
        RECT  5.605 1.640 6.130 1.870 ;
        RECT  5.375 1.190 5.605 1.870 ;
        RECT  4.150 1.190 5.375 1.420 ;
        RECT  4.605 1.655 4.835 2.500 ;
        RECT  3.920 0.990 4.150 2.640 ;
        RECT  3.160 0.465 4.130 0.695 ;
        RECT  3.500 0.990 3.920 1.220 ;
        RECT  3.485 2.410 3.920 2.640 ;
        RECT  2.930 0.465 3.160 1.205 ;
        RECT  2.005 0.975 2.930 1.205 ;
        RECT  1.775 0.975 2.005 2.755 ;
        RECT  1.520 0.975 1.775 1.205 ;
        RECT  1.520 2.525 1.775 2.755 ;
        RECT  1.310 2.985 1.650 3.455 ;
        RECT  0.465 2.985 1.310 3.215 ;
        RECT  0.345 0.980 0.530 1.210 ;
        RECT  0.345 2.425 0.465 3.215 ;
        RECT  0.235 0.980 0.345 3.215 ;
        RECT  0.115 0.980 0.235 2.765 ;
    END
END DFSNQD2BWP7T

MACRO DFXD0BWP7T
    CLASS CORE ;
    FOREIGN DFXD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SA
        ANTENNAGATEAREA 0.5049 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 0.980 2.710 ;
        RECT  0.575 1.730 0.700 2.080 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.075 13.300 2.560 ;
        RECT  12.885 1.075 13.020 1.305 ;
        RECT  12.600 2.330 13.020 2.560 ;
        RECT  12.655 0.520 12.885 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.510 14.420 2.715 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.360 1.605 3.500 1.965 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2250 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.750 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.760 4.900 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.660 0.810 ;
        RECT  10.530 -0.235 13.320 0.235 ;
        RECT  10.190 -0.235 10.530 0.465 ;
        RECT  8.510 -0.235 10.190 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.800 -0.235 4.575 0.235 ;
        RECT  3.460 -0.235 3.800 0.465 ;
        RECT  1.240 -0.235 3.460 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.730 3.685 14.560 4.155 ;
        RECT  13.390 3.365 13.730 4.155 ;
        RECT  11.430 3.685 13.390 4.155 ;
        RECT  11.090 3.385 11.430 4.155 ;
        RECT  8.520 3.685 11.090 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  5.140 3.685 8.160 4.155 ;
        RECT  4.800 3.455 5.140 4.155 ;
        RECT  3.710 3.685 4.800 4.155 ;
        RECT  3.470 2.970 3.710 4.155 ;
        RECT  1.185 3.685 3.470 4.155 ;
        RECT  0.955 2.960 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.020 ;
        RECT  12.370 2.790 13.615 3.020 ;
        RECT  10.990 0.465 12.420 0.695 ;
        RECT  12.140 1.020 12.370 3.020 ;
        RECT  11.450 1.020 12.140 1.250 ;
        RECT  11.900 2.540 12.140 2.775 ;
        RECT  11.680 1.565 11.910 2.310 ;
        RECT  11.450 2.080 11.680 2.310 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  11.220 2.080 11.450 2.995 ;
        RECT  10.735 1.600 11.220 1.830 ;
        RECT  9.935 2.765 11.220 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.500 2.300 10.770 2.530 ;
        RECT  10.500 0.990 10.760 1.220 ;
        RECT  10.270 0.990 10.500 2.530 ;
        RECT  9.225 3.225 10.480 3.455 ;
        RECT  9.705 0.910 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.820 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.590 2.730 7.820 3.455 ;
        RECT  5.845 3.225 7.590 3.455 ;
        RECT  7.035 0.935 7.265 2.915 ;
        RECT  6.315 0.465 6.545 2.830 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  5.845 1.615 6.085 1.955 ;
        RECT  5.615 0.925 5.845 3.455 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.790 ;
        RECT  3.120 0.695 5.145 0.925 ;
        RECT  4.145 1.155 5.140 1.385 ;
        RECT  4.170 2.560 5.140 2.790 ;
        RECT  2.890 0.695 3.120 2.745 ;
        RECT  2.140 0.695 2.890 0.925 ;
        RECT  2.100 2.515 2.890 2.745 ;
        RECT  2.420 1.210 2.650 1.910 ;
        RECT  0.465 1.210 2.420 1.440 ;
        RECT  0.345 0.595 0.465 1.440 ;
        RECT  0.345 2.815 0.465 3.185 ;
        RECT  0.235 0.595 0.345 3.185 ;
        RECT  0.115 1.210 0.235 3.185 ;
    END
END DFXD0BWP7T

MACRO DFXD1BWP7T
    CLASS CORE ;
    FOREIGN DFXD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SA
        ANTENNAGATEAREA 0.5049 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 0.980 2.710 ;
        RECT  0.575 1.730 0.700 2.080 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.075 13.300 2.560 ;
        RECT  12.885 1.075 13.020 1.305 ;
        RECT  12.600 2.330 13.020 2.560 ;
        RECT  12.655 0.480 12.885 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.470 14.420 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.360 1.605 3.500 1.965 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2250 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.750 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.760 4.900 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.660 0.810 ;
        RECT  10.530 -0.235 13.320 0.235 ;
        RECT  10.190 -0.235 10.530 0.465 ;
        RECT  8.510 -0.235 10.190 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.800 -0.235 4.575 0.235 ;
        RECT  3.460 -0.235 3.800 0.465 ;
        RECT  1.240 -0.235 3.460 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 3.685 14.560 4.155 ;
        RECT  13.320 3.250 13.660 4.155 ;
        RECT  11.520 3.685 13.320 4.155 ;
        RECT  11.180 3.250 11.520 4.155 ;
        RECT  8.520 3.685 11.180 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  5.140 3.685 8.160 4.155 ;
        RECT  4.800 3.455 5.140 4.155 ;
        RECT  3.710 3.685 4.800 4.155 ;
        RECT  3.470 2.970 3.710 4.155 ;
        RECT  1.185 3.685 3.470 4.155 ;
        RECT  0.955 2.960 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.020 ;
        RECT  12.370 2.790 13.615 3.020 ;
        RECT  10.990 0.465 12.420 0.695 ;
        RECT  12.185 1.020 12.370 3.020 ;
        RECT  12.140 1.020 12.185 3.380 ;
        RECT  11.450 1.020 12.140 1.250 ;
        RECT  11.955 2.565 12.140 3.380 ;
        RECT  11.680 1.565 11.910 2.310 ;
        RECT  11.450 2.080 11.680 2.310 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  11.220 2.080 11.450 2.995 ;
        RECT  10.735 1.600 11.220 1.830 ;
        RECT  9.935 2.765 11.220 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.500 2.300 10.770 2.530 ;
        RECT  10.500 0.990 10.760 1.220 ;
        RECT  10.270 0.990 10.500 2.530 ;
        RECT  9.225 3.225 10.480 3.455 ;
        RECT  9.705 0.910 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.820 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.590 2.730 7.820 3.455 ;
        RECT  5.845 3.225 7.590 3.455 ;
        RECT  7.035 0.935 7.265 2.915 ;
        RECT  6.315 0.465 6.545 2.830 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  5.845 1.615 6.085 1.955 ;
        RECT  5.615 0.925 5.845 3.455 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.790 ;
        RECT  3.120 0.695 5.145 0.925 ;
        RECT  4.145 1.155 5.140 1.385 ;
        RECT  4.170 2.560 5.140 2.790 ;
        RECT  2.890 0.695 3.120 2.745 ;
        RECT  2.140 0.695 2.890 0.925 ;
        RECT  2.100 2.515 2.890 2.745 ;
        RECT  2.420 1.210 2.650 1.910 ;
        RECT  0.465 1.210 2.420 1.440 ;
        RECT  0.345 0.595 0.465 1.440 ;
        RECT  0.345 2.815 0.465 3.185 ;
        RECT  0.235 0.595 0.345 3.185 ;
        RECT  0.115 1.210 0.235 3.185 ;
    END
END DFXD1BWP7T

MACRO DFXD2BWP7T
    CLASS CORE ;
    FOREIGN DFXD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SA
        ANTENNAGATEAREA 0.5049 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 0.980 2.710 ;
        RECT  0.575 1.730 0.700 2.080 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.560 0.465 13.905 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.055 15.540 2.690 ;
        RECT  15.260 0.465 15.285 3.310 ;
        RECT  15.050 0.465 15.260 1.285 ;
        RECT  15.055 2.460 15.260 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.360 1.605 3.500 1.965 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2250 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.750 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.760 4.900 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.245 ;
        RECT  14.620 -0.235 15.775 0.235 ;
        RECT  14.280 -0.235 14.620 1.180 ;
        RECT  13.140 -0.235 14.280 0.235 ;
        RECT  12.800 -0.235 13.140 0.465 ;
        RECT  11.525 -0.235 12.800 0.235 ;
        RECT  11.185 -0.235 11.525 0.465 ;
        RECT  8.510 -0.235 11.185 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.800 -0.235 4.575 0.235 ;
        RECT  3.460 -0.235 3.800 0.465 ;
        RECT  1.240 -0.235 3.460 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.255 16.005 4.155 ;
        RECT  14.620 3.685 15.775 4.155 ;
        RECT  14.280 3.250 14.620 4.155 ;
        RECT  13.105 3.685 14.280 4.155 ;
        RECT  12.765 3.250 13.105 4.155 ;
        RECT  11.575 3.685 12.765 4.155 ;
        RECT  11.235 3.250 11.575 4.155 ;
        RECT  8.520 3.685 11.235 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  5.140 3.685 8.160 4.155 ;
        RECT  4.800 3.455 5.140 4.155 ;
        RECT  3.710 3.685 4.800 4.155 ;
        RECT  3.470 2.970 3.710 4.155 ;
        RECT  1.185 3.685 3.470 4.155 ;
        RECT  0.955 2.960 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.575 1.600 14.805 3.010 ;
        RECT  12.555 2.780 14.575 3.010 ;
        RECT  13.090 0.695 13.320 1.940 ;
        RECT  10.990 0.695 13.090 0.925 ;
        RECT  12.325 1.155 12.555 3.010 ;
        RECT  11.505 1.155 12.325 1.385 ;
        RECT  12.285 2.565 12.325 3.010 ;
        RECT  12.055 2.565 12.285 3.380 ;
        RECT  11.800 1.675 12.030 2.310 ;
        RECT  11.530 2.080 11.800 2.310 ;
        RECT  11.300 2.080 11.530 2.995 ;
        RECT  11.275 1.155 11.505 1.830 ;
        RECT  9.935 2.765 11.300 2.995 ;
        RECT  10.725 1.600 11.275 1.830 ;
        RECT  10.760 0.695 10.990 1.220 ;
        RECT  10.460 2.300 10.770 2.530 ;
        RECT  10.460 0.990 10.760 1.220 ;
        RECT  10.230 0.990 10.460 2.530 ;
        RECT  9.225 3.225 10.425 3.455 ;
        RECT  9.705 0.935 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.820 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.590 2.730 7.820 3.455 ;
        RECT  5.845 3.225 7.590 3.455 ;
        RECT  7.035 0.935 7.265 2.915 ;
        RECT  6.315 0.465 6.545 2.830 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  5.845 1.615 6.085 1.955 ;
        RECT  5.615 0.925 5.845 3.455 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.790 ;
        RECT  3.120 0.695 5.145 0.925 ;
        RECT  4.145 1.155 5.140 1.385 ;
        RECT  4.170 2.560 5.140 2.790 ;
        RECT  2.890 0.695 3.120 2.745 ;
        RECT  2.140 0.695 2.890 0.925 ;
        RECT  2.100 2.515 2.890 2.745 ;
        RECT  2.420 1.210 2.650 1.910 ;
        RECT  0.465 1.210 2.420 1.440 ;
        RECT  0.345 0.595 0.465 1.440 ;
        RECT  0.345 2.815 0.465 3.185 ;
        RECT  0.235 0.595 0.345 3.185 ;
        RECT  0.115 1.210 0.235 3.185 ;
    END
END DFXD2BWP7T

MACRO DFXQD1BWP7T
    CLASS CORE ;
    FOREIGN DFXQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SA
        ANTENNAGATEAREA 0.5049 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 0.980 2.710 ;
        RECT  0.575 1.730 0.700 2.080 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.530 0.470 13.860 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.370 1.605 3.500 1.965 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2637 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.725 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.760 4.910 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.050 -0.235 14.000 0.235 ;
        RECT  12.810 -0.235 13.050 1.260 ;
        RECT  11.635 -0.235 12.810 0.235 ;
        RECT  11.295 -0.235 11.635 0.780 ;
        RECT  8.595 -0.235 11.295 0.235 ;
        RECT  8.255 -0.235 8.595 0.730 ;
        RECT  4.925 -0.235 8.255 0.235 ;
        RECT  4.585 -0.235 4.925 0.465 ;
        RECT  3.810 -0.235 4.585 0.235 ;
        RECT  3.470 -0.235 3.810 0.465 ;
        RECT  1.240 -0.235 3.470 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.045 3.685 14.000 4.155 ;
        RECT  12.815 2.250 13.045 4.155 ;
        RECT  11.635 3.685 12.815 4.155 ;
        RECT  11.295 3.250 11.635 4.155 ;
        RECT  8.605 3.685 11.295 4.155 ;
        RECT  8.245 3.190 8.605 4.155 ;
        RECT  5.150 3.685 8.245 4.155 ;
        RECT  4.810 3.455 5.150 4.155 ;
        RECT  3.720 3.685 4.810 4.155 ;
        RECT  3.480 2.950 3.720 4.155 ;
        RECT  1.185 3.685 3.480 4.155 ;
        RECT  0.955 2.960 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.530 1.600 13.285 1.945 ;
        RECT  12.350 1.020 12.530 2.825 ;
        RECT  12.345 0.490 12.350 2.825 ;
        RECT  12.300 0.490 12.345 3.380 ;
        RECT  12.115 0.490 12.300 1.250 ;
        RECT  12.115 2.565 12.300 3.380 ;
        RECT  11.450 1.020 12.115 1.250 ;
        RECT  11.840 1.605 12.070 2.310 ;
        RECT  11.565 2.080 11.840 2.310 ;
        RECT  11.335 2.080 11.565 2.995 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  10.050 2.765 11.335 2.995 ;
        RECT  10.850 1.600 11.220 1.830 ;
        RECT  10.615 2.300 10.885 2.530 ;
        RECT  10.615 0.990 10.835 1.220 ;
        RECT  10.385 0.990 10.615 2.530 ;
        RECT  9.340 3.225 10.595 3.455 ;
        RECT  9.820 0.910 10.050 2.995 ;
        RECT  9.360 0.960 9.590 2.500 ;
        RECT  8.260 0.960 9.360 1.190 ;
        RECT  9.045 2.270 9.360 2.500 ;
        RECT  9.110 2.730 9.340 3.455 ;
        RECT  7.855 2.730 9.110 2.960 ;
        RECT  8.785 1.560 9.090 1.900 ;
        RECT  8.555 1.560 8.785 2.415 ;
        RECT  7.300 2.185 8.555 2.415 ;
        RECT  8.030 0.960 8.260 1.890 ;
        RECT  7.625 2.730 7.855 3.415 ;
        RECT  5.880 3.185 7.625 3.415 ;
        RECT  7.070 0.935 7.300 2.915 ;
        RECT  6.350 0.465 6.580 2.830 ;
        RECT  5.385 0.465 6.350 0.695 ;
        RECT  5.880 1.615 6.120 1.955 ;
        RECT  5.650 0.925 5.880 3.415 ;
        RECT  5.155 0.465 5.385 0.925 ;
        RECT  5.150 1.155 5.380 2.790 ;
        RECT  3.130 0.695 5.155 0.925 ;
        RECT  4.155 1.155 5.150 1.385 ;
        RECT  4.180 2.560 5.150 2.790 ;
        RECT  2.900 0.695 3.130 2.745 ;
        RECT  2.150 0.695 2.900 0.925 ;
        RECT  2.110 2.515 2.900 2.745 ;
        RECT  2.430 1.210 2.660 1.910 ;
        RECT  0.465 1.210 2.430 1.440 ;
        RECT  0.345 0.595 0.465 1.440 ;
        RECT  0.345 2.815 0.465 3.185 ;
        RECT  0.235 0.595 0.345 3.185 ;
        RECT  0.115 1.210 0.235 3.185 ;
    END
END DFXQD1BWP7T

MACRO DFXQD2BWP7T
    CLASS CORE ;
    FOREIGN DFXQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SA
        ANTENNAGATEAREA 0.5049 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 0.980 2.710 ;
        RECT  0.575 1.730 0.700 2.080 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.605 1.060 13.860 2.715 ;
        RECT  13.580 0.480 13.605 3.310 ;
        RECT  13.375 0.480 13.580 1.290 ;
        RECT  13.375 2.480 13.580 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.370 1.605 3.500 1.965 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2637 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.725 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.760 4.910 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 -0.235 14.560 0.235 ;
        RECT  14.095 -0.235 14.325 1.240 ;
        RECT  12.900 -0.235 14.095 0.235 ;
        RECT  12.560 -0.235 12.900 0.465 ;
        RECT  11.585 -0.235 12.560 0.235 ;
        RECT  11.245 -0.235 11.585 0.780 ;
        RECT  8.595 -0.235 11.245 0.235 ;
        RECT  8.255 -0.235 8.595 0.730 ;
        RECT  4.925 -0.235 8.255 0.235 ;
        RECT  4.585 -0.235 4.925 0.465 ;
        RECT  3.810 -0.235 4.585 0.235 ;
        RECT  3.470 -0.235 3.810 0.465 ;
        RECT  1.240 -0.235 3.470 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 3.685 14.560 4.155 ;
        RECT  14.095 2.255 14.325 4.155 ;
        RECT  12.940 3.685 14.095 4.155 ;
        RECT  12.600 3.240 12.940 4.155 ;
        RECT  11.635 3.685 12.600 4.155 ;
        RECT  11.295 3.250 11.635 4.155 ;
        RECT  8.605 3.685 11.295 4.155 ;
        RECT  8.245 3.190 8.605 4.155 ;
        RECT  5.150 3.685 8.245 4.155 ;
        RECT  4.810 3.455 5.150 4.155 ;
        RECT  3.720 3.685 4.810 4.155 ;
        RECT  3.480 2.950 3.720 4.155 ;
        RECT  1.185 3.685 3.480 4.155 ;
        RECT  0.955 2.960 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.730 1.600 13.125 1.945 ;
        RECT  12.500 1.020 12.730 2.795 ;
        RECT  11.450 1.020 12.500 1.250 ;
        RECT  12.015 2.565 12.500 2.795 ;
        RECT  11.840 1.605 12.070 2.310 ;
        RECT  11.565 2.080 11.840 2.310 ;
        RECT  11.335 2.080 11.565 2.995 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  10.050 2.765 11.335 2.995 ;
        RECT  10.850 1.600 11.220 1.830 ;
        RECT  10.615 2.300 10.885 2.530 ;
        RECT  10.615 0.990 10.835 1.220 ;
        RECT  10.385 0.990 10.615 2.530 ;
        RECT  9.340 3.225 10.595 3.455 ;
        RECT  9.820 0.910 10.050 2.995 ;
        RECT  9.360 0.960 9.590 2.500 ;
        RECT  8.260 0.960 9.360 1.190 ;
        RECT  9.045 2.270 9.360 2.500 ;
        RECT  9.110 2.730 9.340 3.455 ;
        RECT  7.855 2.730 9.110 2.960 ;
        RECT  8.785 1.560 9.090 1.900 ;
        RECT  8.555 1.560 8.785 2.415 ;
        RECT  7.300 2.185 8.555 2.415 ;
        RECT  8.030 0.960 8.260 1.890 ;
        RECT  7.625 2.730 7.855 3.415 ;
        RECT  5.880 3.185 7.625 3.415 ;
        RECT  7.070 0.935 7.300 2.915 ;
        RECT  6.350 0.465 6.580 2.830 ;
        RECT  5.385 0.465 6.350 0.695 ;
        RECT  5.880 1.615 6.120 1.955 ;
        RECT  5.650 0.925 5.880 3.415 ;
        RECT  5.155 0.465 5.385 0.925 ;
        RECT  5.150 1.155 5.380 2.790 ;
        RECT  3.130 0.695 5.155 0.925 ;
        RECT  4.155 1.155 5.150 1.385 ;
        RECT  4.180 2.560 5.150 2.790 ;
        RECT  2.900 0.695 3.130 2.745 ;
        RECT  2.150 0.695 2.900 0.925 ;
        RECT  2.110 2.515 2.900 2.745 ;
        RECT  2.430 1.210 2.660 1.910 ;
        RECT  0.465 1.210 2.430 1.440 ;
        RECT  0.345 0.595 0.465 1.440 ;
        RECT  0.345 2.815 0.465 3.185 ;
        RECT  0.235 0.595 0.345 3.185 ;
        RECT  0.115 1.210 0.235 3.185 ;
    END
END DFXQD2BWP7T

MACRO EDFCND0BWP7T
    CLASS CORE ;
    FOREIGN EDFCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.075 15.540 2.560 ;
        RECT  15.125 1.075 15.260 1.305 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.545 15.125 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.515 16.660 2.775 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.3942 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.240 2.395 13.355 2.625 ;
        RECT  13.010 2.395 13.240 3.455 ;
        RECT  10.830 3.225 13.010 3.455 ;
        RECT  10.600 2.730 10.830 3.455 ;
        RECT  9.670 2.730 10.600 2.960 ;
        RECT  9.440 2.730 9.670 3.270 ;
        RECT  7.665 2.940 9.440 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.810 ;
        RECT  12.125 -0.235 15.560 0.235 ;
        RECT  11.785 -0.235 12.125 0.465 ;
        RECT  8.695 -0.235 11.785 0.235 ;
        RECT  8.355 -0.235 8.695 0.730 ;
        RECT  4.550 -0.235 8.355 0.235 ;
        RECT  4.210 -0.235 4.550 0.465 ;
        RECT  3.660 -0.235 4.210 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 3.685 16.800 4.155 ;
        RECT  15.560 3.305 15.900 4.155 ;
        RECT  14.640 3.685 15.560 4.155 ;
        RECT  14.300 3.455 14.640 4.155 ;
        RECT  10.360 3.685 14.300 4.155 ;
        RECT  10.020 3.190 10.360 4.155 ;
        RECT  3.945 3.685 10.020 4.155 ;
        RECT  3.605 3.440 3.945 4.155 ;
        RECT  1.250 3.685 3.605 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  14.575 2.790 15.855 3.020 ;
        RECT  12.805 0.465 14.660 0.695 ;
        RECT  14.345 1.020 14.575 3.020 ;
        RECT  13.490 1.020 14.345 1.250 ;
        RECT  13.820 2.390 14.345 2.620 ;
        RECT  13.835 1.565 14.065 2.160 ;
        RECT  12.735 1.930 13.835 2.160 ;
        RECT  13.590 2.390 13.820 3.200 ;
        RECT  13.260 1.020 13.490 1.700 ;
        RECT  12.235 1.470 13.260 1.700 ;
        RECT  12.575 0.465 12.805 1.180 ;
        RECT  12.505 1.930 12.735 2.995 ;
        RECT  11.955 0.950 12.575 1.180 ;
        RECT  11.295 2.765 12.505 2.995 ;
        RECT  11.955 2.305 12.225 2.535 ;
        RECT  11.725 0.950 11.955 2.535 ;
        RECT  11.045 0.950 11.725 1.220 ;
        RECT  11.065 1.615 11.295 2.995 ;
        RECT  10.490 1.615 11.065 1.845 ;
        RECT  10.815 0.465 11.045 1.220 ;
        RECT  9.155 0.465 10.815 0.695 ;
        RECT  10.260 0.990 10.490 1.845 ;
        RECT  9.870 2.270 10.385 2.500 ;
        RECT  10.030 0.990 10.260 1.220 ;
        RECT  9.640 1.420 9.870 2.500 ;
        RECT  9.615 1.420 9.640 1.650 ;
        RECT  9.385 0.925 9.615 1.650 ;
        RECT  8.605 1.420 9.385 1.650 ;
        RECT  8.935 1.880 9.275 2.200 ;
        RECT  8.925 0.465 9.155 1.190 ;
        RECT  7.425 2.440 9.085 2.670 ;
        RECT  6.905 1.970 8.935 2.200 ;
        RECT  7.660 0.960 8.925 1.190 ;
        RECT  8.265 1.420 8.605 1.740 ;
        RECT  7.430 0.465 7.660 1.190 ;
        RECT  5.015 0.465 7.430 0.695 ;
        RECT  6.900 1.970 6.905 2.725 ;
        RECT  6.670 0.935 6.900 2.725 ;
        RECT  6.135 0.925 6.270 2.865 ;
        RECT  6.035 0.925 6.135 3.210 ;
        RECT  5.845 0.925 6.035 1.155 ;
        RECT  5.905 2.525 6.035 3.210 ;
        RECT  2.675 2.980 5.905 3.210 ;
        RECT  5.605 1.805 5.805 2.035 ;
        RECT  5.375 1.115 5.605 2.715 ;
        RECT  5.145 1.115 5.375 1.345 ;
        RECT  5.150 2.485 5.375 2.715 ;
        RECT  4.885 1.800 5.080 2.040 ;
        RECT  4.785 0.465 5.015 0.925 ;
        RECT  4.655 1.155 4.885 2.670 ;
        RECT  3.175 0.695 4.785 0.925 ;
        RECT  3.820 1.155 4.655 1.385 ;
        RECT  3.790 2.435 4.655 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.745 2.675 3.210 ;
        RECT  2.060 0.745 2.445 0.975 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFCND0BWP7T

MACRO EDFCND1BWP7T
    CLASS CORE ;
    FOREIGN EDFCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.9672 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.075 15.540 2.560 ;
        RECT  15.125 1.075 15.260 1.305 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.480 15.125 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.470 16.660 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.3942 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.240 2.395 13.355 2.625 ;
        RECT  13.010 2.395 13.240 3.455 ;
        RECT  10.830 3.225 13.010 3.455 ;
        RECT  10.600 2.730 10.830 3.455 ;
        RECT  9.670 2.730 10.600 2.960 ;
        RECT  9.440 2.730 9.670 3.270 ;
        RECT  7.665 2.940 9.440 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.810 ;
        RECT  12.125 -0.235 15.560 0.235 ;
        RECT  11.785 -0.235 12.125 0.465 ;
        RECT  8.695 -0.235 11.785 0.235 ;
        RECT  8.355 -0.235 8.695 0.730 ;
        RECT  4.550 -0.235 8.355 0.235 ;
        RECT  4.210 -0.235 4.550 0.465 ;
        RECT  3.660 -0.235 4.210 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 3.685 16.800 4.155 ;
        RECT  15.560 3.250 15.900 4.155 ;
        RECT  14.640 3.685 15.560 4.155 ;
        RECT  14.300 3.455 14.640 4.155 ;
        RECT  10.360 3.685 14.300 4.155 ;
        RECT  10.020 3.190 10.360 4.155 ;
        RECT  3.945 3.685 10.020 4.155 ;
        RECT  3.605 3.440 3.945 4.155 ;
        RECT  1.250 3.685 3.605 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  14.575 2.790 15.855 3.020 ;
        RECT  12.805 0.465 14.660 0.695 ;
        RECT  14.345 1.020 14.575 3.020 ;
        RECT  13.490 1.020 14.345 1.250 ;
        RECT  13.820 2.390 14.345 2.620 ;
        RECT  13.835 1.565 14.065 2.160 ;
        RECT  12.735 1.930 13.835 2.160 ;
        RECT  13.590 2.390 13.820 3.200 ;
        RECT  13.260 1.020 13.490 1.700 ;
        RECT  12.235 1.470 13.260 1.700 ;
        RECT  12.575 0.465 12.805 1.180 ;
        RECT  12.505 1.930 12.735 2.995 ;
        RECT  11.955 0.950 12.575 1.180 ;
        RECT  11.295 2.765 12.505 2.995 ;
        RECT  11.955 2.305 12.225 2.535 ;
        RECT  11.725 0.950 11.955 2.535 ;
        RECT  11.045 0.950 11.725 1.220 ;
        RECT  11.065 1.615 11.295 2.995 ;
        RECT  10.490 1.615 11.065 1.845 ;
        RECT  10.815 0.465 11.045 1.220 ;
        RECT  9.155 0.465 10.815 0.695 ;
        RECT  10.260 0.990 10.490 1.845 ;
        RECT  9.870 2.270 10.385 2.500 ;
        RECT  10.030 0.990 10.260 1.220 ;
        RECT  9.640 1.420 9.870 2.500 ;
        RECT  9.615 1.420 9.640 1.650 ;
        RECT  9.385 0.925 9.615 1.650 ;
        RECT  8.605 1.420 9.385 1.650 ;
        RECT  8.935 1.880 9.275 2.200 ;
        RECT  8.925 0.465 9.155 1.190 ;
        RECT  7.425 2.440 9.085 2.670 ;
        RECT  6.905 1.970 8.935 2.200 ;
        RECT  7.660 0.960 8.925 1.190 ;
        RECT  8.265 1.420 8.605 1.740 ;
        RECT  7.430 0.465 7.660 1.190 ;
        RECT  5.015 0.465 7.430 0.695 ;
        RECT  6.900 1.970 6.905 2.725 ;
        RECT  6.670 0.935 6.900 2.725 ;
        RECT  6.135 0.925 6.270 2.865 ;
        RECT  6.035 0.925 6.135 3.210 ;
        RECT  5.845 0.925 6.035 1.155 ;
        RECT  5.905 2.525 6.035 3.210 ;
        RECT  2.675 2.980 5.905 3.210 ;
        RECT  5.605 1.805 5.805 2.035 ;
        RECT  5.375 1.115 5.605 2.715 ;
        RECT  5.145 1.115 5.375 1.345 ;
        RECT  5.150 2.485 5.375 2.715 ;
        RECT  4.885 1.800 5.080 2.040 ;
        RECT  4.785 0.465 5.015 0.925 ;
        RECT  4.655 1.155 4.885 2.670 ;
        RECT  3.175 0.695 4.785 0.925 ;
        RECT  3.820 1.155 4.655 1.385 ;
        RECT  3.790 2.435 4.655 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.745 2.675 3.210 ;
        RECT  2.060 0.745 2.445 0.975 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFCND1BWP7T

MACRO EDFCND2BWP7T
    CLASS CORE ;
    FOREIGN EDFCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.100 2.235 16.140 2.560 ;
        RECT  15.820 0.480 16.100 2.560 ;
        RECT  15.800 2.245 15.820 2.560 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.525 1.075 17.780 2.715 ;
        RECT  17.500 0.480 17.525 3.455 ;
        RECT  17.295 0.480 17.500 1.305 ;
        RECT  17.295 2.445 17.500 3.455 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.3942 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.990 3.085 13.335 3.455 ;
        RECT  10.830 3.225 12.990 3.455 ;
        RECT  10.600 2.730 10.830 3.455 ;
        RECT  9.670 2.730 10.600 2.960 ;
        RECT  9.440 2.730 9.670 3.270 ;
        RECT  7.665 2.940 9.440 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 -0.235 18.480 0.235 ;
        RECT  18.015 -0.235 18.245 1.300 ;
        RECT  16.805 -0.235 18.015 0.235 ;
        RECT  16.575 -0.235 16.805 1.290 ;
        RECT  15.365 -0.235 16.575 0.235 ;
        RECT  15.135 -0.235 15.365 0.780 ;
        RECT  12.735 -0.235 15.135 0.235 ;
        RECT  12.505 -0.235 12.735 0.725 ;
        RECT  8.695 -0.235 12.505 0.235 ;
        RECT  8.355 -0.235 8.695 0.730 ;
        RECT  4.550 -0.235 8.355 0.235 ;
        RECT  4.210 -0.235 4.550 0.465 ;
        RECT  3.660 -0.235 4.210 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 3.685 18.480 4.155 ;
        RECT  18.015 2.245 18.245 4.155 ;
        RECT  16.860 3.685 18.015 4.155 ;
        RECT  16.520 3.250 16.860 4.155 ;
        RECT  15.420 3.685 16.520 4.155 ;
        RECT  15.080 3.250 15.420 4.155 ;
        RECT  13.965 3.685 15.080 4.155 ;
        RECT  13.625 3.455 13.965 4.155 ;
        RECT  10.360 3.685 13.625 4.155 ;
        RECT  10.020 3.190 10.360 4.155 ;
        RECT  3.945 3.685 10.020 4.155 ;
        RECT  3.605 3.440 3.945 4.155 ;
        RECT  1.250 3.685 3.605 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.815 1.600 17.045 3.020 ;
        RECT  15.395 2.790 16.815 3.020 ;
        RECT  15.165 1.020 15.395 3.020 ;
        RECT  13.795 1.020 15.165 1.250 ;
        RECT  14.645 2.445 15.165 2.675 ;
        RECT  13.335 0.560 14.905 0.790 ;
        RECT  14.415 2.445 14.645 3.380 ;
        RECT  13.485 2.445 14.415 2.675 ;
        RECT  14.115 1.640 14.345 2.160 ;
        RECT  12.735 1.930 14.115 2.160 ;
        RECT  13.565 1.020 13.795 1.645 ;
        RECT  12.245 1.415 13.565 1.645 ;
        RECT  13.105 0.560 13.335 1.185 ;
        RECT  11.755 0.955 13.105 1.185 ;
        RECT  12.505 1.930 12.735 2.995 ;
        RECT  11.295 2.765 12.505 2.995 ;
        RECT  12.015 1.415 12.245 1.940 ;
        RECT  11.755 2.300 12.070 2.530 ;
        RECT  11.525 0.955 11.755 2.530 ;
        RECT  11.110 0.955 11.525 1.220 ;
        RECT  11.065 1.615 11.295 2.995 ;
        RECT  10.815 0.465 11.110 1.220 ;
        RECT  10.490 1.615 11.065 1.845 ;
        RECT  9.155 0.465 10.815 0.695 ;
        RECT  10.260 0.990 10.490 1.845 ;
        RECT  9.870 2.270 10.385 2.500 ;
        RECT  10.030 0.990 10.260 1.220 ;
        RECT  9.640 1.420 9.870 2.500 ;
        RECT  9.615 1.420 9.640 1.650 ;
        RECT  9.385 0.925 9.615 1.650 ;
        RECT  8.605 1.420 9.385 1.650 ;
        RECT  8.935 1.880 9.275 2.200 ;
        RECT  8.925 0.465 9.155 1.190 ;
        RECT  7.425 2.440 9.085 2.670 ;
        RECT  6.905 1.970 8.935 2.200 ;
        RECT  7.660 0.960 8.925 1.190 ;
        RECT  8.265 1.420 8.605 1.740 ;
        RECT  7.430 0.465 7.660 1.190 ;
        RECT  5.015 0.465 7.430 0.695 ;
        RECT  6.900 1.970 6.905 2.725 ;
        RECT  6.670 0.935 6.900 2.725 ;
        RECT  6.135 0.925 6.270 2.865 ;
        RECT  6.035 0.925 6.135 3.210 ;
        RECT  5.845 0.925 6.035 1.155 ;
        RECT  5.905 2.525 6.035 3.210 ;
        RECT  2.675 2.980 5.905 3.210 ;
        RECT  5.605 1.805 5.805 2.035 ;
        RECT  5.375 1.115 5.605 2.715 ;
        RECT  5.145 1.115 5.375 1.345 ;
        RECT  5.150 2.485 5.375 2.715 ;
        RECT  4.885 1.800 5.080 2.040 ;
        RECT  4.785 0.465 5.015 0.925 ;
        RECT  4.655 1.155 4.885 2.670 ;
        RECT  3.175 0.695 4.785 0.925 ;
        RECT  3.820 1.155 4.655 1.385 ;
        RECT  3.790 2.435 4.655 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.745 2.675 3.210 ;
        RECT  2.060 0.745 2.445 0.975 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFCND2BWP7T

MACRO EDFCNQD1BWP7T
    CLASS CORE ;
    FOREIGN EDFCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.210 0.470 15.540 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.3942 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.130 2.395 13.245 2.625 ;
        RECT  12.900 2.395 13.130 3.455 ;
        RECT  10.830 3.225 12.900 3.455 ;
        RECT  10.600 2.730 10.830 3.455 ;
        RECT  9.670 2.730 10.600 2.960 ;
        RECT  9.440 2.730 9.670 3.270 ;
        RECT  7.665 2.940 9.440 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.780 -0.235 15.680 0.235 ;
        RECT  14.440 -0.235 14.780 0.790 ;
        RECT  12.755 -0.235 14.440 0.235 ;
        RECT  12.415 -0.235 12.755 1.180 ;
        RECT  8.695 -0.235 12.415 0.235 ;
        RECT  8.355 -0.235 8.695 0.730 ;
        RECT  4.550 -0.235 8.355 0.235 ;
        RECT  4.210 -0.235 4.550 0.465 ;
        RECT  3.660 -0.235 4.210 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.585 3.685 15.680 4.155 ;
        RECT  14.240 2.900 14.585 4.155 ;
        RECT  10.360 3.685 14.240 4.155 ;
        RECT  10.020 3.190 10.360 4.155 ;
        RECT  3.945 3.685 10.020 4.155 ;
        RECT  3.605 3.440 3.945 4.155 ;
        RECT  1.250 3.685 3.605 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.465 1.600 14.965 1.940 ;
        RECT  14.235 1.020 14.465 2.620 ;
        RECT  14.080 1.020 14.235 1.250 ;
        RECT  13.710 2.390 14.235 2.620 ;
        RECT  13.720 0.545 14.080 1.250 ;
        RECT  13.725 1.565 13.955 2.160 ;
        RECT  12.670 1.930 13.725 2.160 ;
        RECT  13.325 1.020 13.720 1.250 ;
        RECT  13.480 2.390 13.710 3.200 ;
        RECT  13.095 1.020 13.325 1.700 ;
        RECT  12.170 1.470 13.095 1.700 ;
        RECT  12.440 1.930 12.670 2.995 ;
        RECT  11.295 2.765 12.440 2.995 ;
        RECT  11.890 2.305 12.160 2.535 ;
        RECT  11.890 0.950 11.975 1.180 ;
        RECT  11.660 0.950 11.890 2.535 ;
        RECT  11.045 0.950 11.660 1.220 ;
        RECT  11.065 1.615 11.295 2.995 ;
        RECT  10.490 1.615 11.065 1.845 ;
        RECT  10.815 0.465 11.045 1.220 ;
        RECT  9.155 0.465 10.815 0.695 ;
        RECT  10.260 0.990 10.490 1.845 ;
        RECT  9.870 2.270 10.385 2.500 ;
        RECT  10.030 0.990 10.260 1.220 ;
        RECT  9.640 1.420 9.870 2.500 ;
        RECT  9.615 1.420 9.640 1.650 ;
        RECT  9.385 0.925 9.615 1.650 ;
        RECT  8.605 1.420 9.385 1.650 ;
        RECT  8.935 1.880 9.275 2.200 ;
        RECT  8.925 0.465 9.155 1.190 ;
        RECT  7.425 2.440 9.085 2.670 ;
        RECT  6.905 1.970 8.935 2.200 ;
        RECT  7.660 0.960 8.925 1.190 ;
        RECT  8.265 1.420 8.605 1.740 ;
        RECT  7.430 0.465 7.660 1.190 ;
        RECT  5.015 0.465 7.430 0.695 ;
        RECT  6.900 1.970 6.905 2.725 ;
        RECT  6.670 0.935 6.900 2.725 ;
        RECT  6.135 0.925 6.270 2.865 ;
        RECT  6.035 0.925 6.135 3.210 ;
        RECT  5.845 0.925 6.035 1.155 ;
        RECT  5.905 2.525 6.035 3.210 ;
        RECT  2.675 2.980 5.905 3.210 ;
        RECT  5.605 1.805 5.805 2.035 ;
        RECT  5.375 1.115 5.605 2.715 ;
        RECT  5.145 1.115 5.375 1.345 ;
        RECT  5.150 2.485 5.375 2.715 ;
        RECT  4.885 1.800 5.080 2.040 ;
        RECT  4.785 0.465 5.015 0.925 ;
        RECT  4.655 1.155 4.885 2.670 ;
        RECT  3.175 0.695 4.785 0.925 ;
        RECT  3.820 1.155 4.655 1.385 ;
        RECT  3.790 2.435 4.655 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.745 2.675 3.210 ;
        RECT  2.060 0.745 2.445 0.975 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFCNQD1BWP7T

MACRO EDFCNQD2BWP7T
    CLASS CORE ;
    FOREIGN EDFCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.845 1.065 16.100 2.620 ;
        RECT  15.820 0.480 15.845 3.310 ;
        RECT  15.615 0.480 15.820 1.360 ;
        RECT  15.615 2.325 15.820 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.3942 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.900 3.085 13.245 3.455 ;
        RECT  10.830 3.225 12.900 3.455 ;
        RECT  10.600 2.730 10.830 3.455 ;
        RECT  9.670 2.730 10.600 2.960 ;
        RECT  9.440 2.730 9.670 3.270 ;
        RECT  7.665 2.940 9.440 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.565 -0.235 16.800 0.235 ;
        RECT  16.335 -0.235 16.565 1.300 ;
        RECT  15.125 -0.235 16.335 0.235 ;
        RECT  14.895 -0.235 15.125 1.300 ;
        RECT  12.700 -0.235 14.895 0.235 ;
        RECT  12.470 -0.235 12.700 1.235 ;
        RECT  8.695 -0.235 12.470 0.235 ;
        RECT  8.355 -0.235 8.695 0.730 ;
        RECT  4.550 -0.235 8.355 0.235 ;
        RECT  4.210 -0.235 4.550 0.465 ;
        RECT  3.660 -0.235 4.210 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.565 3.685 16.800 4.155 ;
        RECT  16.335 2.235 16.565 4.155 ;
        RECT  15.125 3.685 16.335 4.155 ;
        RECT  14.895 2.245 15.125 4.155 ;
        RECT  13.705 3.685 14.895 4.155 ;
        RECT  13.475 3.400 13.705 4.155 ;
        RECT  10.360 3.685 13.475 4.155 ;
        RECT  10.020 3.190 10.360 4.155 ;
        RECT  3.945 3.685 10.020 4.155 ;
        RECT  3.605 3.440 3.945 4.155 ;
        RECT  1.250 3.685 3.605 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.425 1.600 15.585 1.940 ;
        RECT  14.405 1.020 14.425 1.940 ;
        RECT  14.175 1.020 14.405 3.395 ;
        RECT  14.170 1.020 14.175 1.250 ;
        RECT  13.120 2.565 14.175 2.795 ;
        RECT  13.940 0.495 14.170 1.250 ;
        RECT  13.715 1.565 13.945 2.310 ;
        RECT  13.160 1.020 13.940 1.250 ;
        RECT  12.670 2.080 13.715 2.310 ;
        RECT  12.930 1.020 13.160 1.850 ;
        RECT  12.225 1.510 12.930 1.850 ;
        RECT  12.440 2.080 12.670 2.995 ;
        RECT  11.295 2.765 12.440 2.995 ;
        RECT  11.975 2.300 12.070 2.530 ;
        RECT  11.730 0.950 11.975 2.530 ;
        RECT  11.045 0.950 11.730 1.220 ;
        RECT  11.065 1.615 11.295 2.995 ;
        RECT  10.490 1.615 11.065 1.845 ;
        RECT  10.815 0.465 11.045 1.220 ;
        RECT  9.155 0.465 10.815 0.695 ;
        RECT  10.260 0.990 10.490 1.845 ;
        RECT  9.870 2.270 10.385 2.500 ;
        RECT  10.030 0.990 10.260 1.220 ;
        RECT  9.640 1.420 9.870 2.500 ;
        RECT  9.615 1.420 9.640 1.650 ;
        RECT  9.385 0.925 9.615 1.650 ;
        RECT  8.605 1.420 9.385 1.650 ;
        RECT  8.935 1.880 9.275 2.200 ;
        RECT  8.925 0.465 9.155 1.190 ;
        RECT  7.425 2.440 9.085 2.670 ;
        RECT  6.905 1.970 8.935 2.200 ;
        RECT  7.660 0.960 8.925 1.190 ;
        RECT  8.265 1.420 8.605 1.740 ;
        RECT  7.430 0.465 7.660 1.190 ;
        RECT  5.015 0.465 7.430 0.695 ;
        RECT  6.900 1.970 6.905 2.725 ;
        RECT  6.670 0.935 6.900 2.725 ;
        RECT  6.135 0.925 6.270 2.865 ;
        RECT  6.035 0.925 6.135 3.210 ;
        RECT  5.845 0.925 6.035 1.155 ;
        RECT  5.905 2.525 6.035 3.210 ;
        RECT  2.675 2.980 5.905 3.210 ;
        RECT  5.605 1.805 5.805 2.035 ;
        RECT  5.375 1.115 5.605 2.715 ;
        RECT  5.145 1.115 5.375 1.345 ;
        RECT  5.150 2.485 5.375 2.715 ;
        RECT  4.885 1.800 5.080 2.040 ;
        RECT  4.785 0.465 5.015 0.925 ;
        RECT  4.655 1.155 4.885 2.670 ;
        RECT  3.175 0.695 4.785 0.925 ;
        RECT  3.820 1.155 4.655 1.385 ;
        RECT  3.790 2.435 4.655 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.745 2.675 3.210 ;
        RECT  2.060 0.745 2.445 0.975 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFCNQD2BWP7T

MACRO EDFD0BWP7T
    CLASS CORE ;
    FOREIGN EDFD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5608 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.475 13.300 2.730 ;
        RECT  12.885 1.475 13.020 1.705 ;
        RECT  12.600 2.500 13.020 2.730 ;
        RECT  12.655 0.920 12.885 1.705 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.940 14.420 2.770 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.605 -0.235 14.560 0.235 ;
        RECT  13.375 -0.235 13.605 1.225 ;
        RECT  10.530 -0.235 13.375 0.235 ;
        RECT  10.300 -0.235 10.530 0.520 ;
        RECT  7.945 -0.235 10.300 0.235 ;
        RECT  7.715 -0.235 7.945 0.785 ;
        RECT  4.360 -0.235 7.715 0.235 ;
        RECT  4.020 -0.235 4.360 0.465 ;
        RECT  3.660 -0.235 4.020 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.700 3.685 14.560 4.155 ;
        RECT  13.360 3.420 13.700 4.155 ;
        RECT  11.515 3.685 13.360 4.155 ;
        RECT  11.170 3.300 11.515 4.155 ;
        RECT  8.185 3.685 11.170 4.155 ;
        RECT  7.825 3.190 8.185 4.155 ;
        RECT  4.680 3.685 7.825 4.155 ;
        RECT  4.340 3.455 4.680 4.155 ;
        RECT  3.620 3.685 4.340 4.155 ;
        RECT  3.280 3.455 3.620 4.155 ;
        RECT  1.250 3.685 3.280 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.190 ;
        RECT  12.370 2.960 13.615 3.190 ;
        RECT  10.990 0.465 12.580 0.695 ;
        RECT  12.140 0.990 12.370 3.190 ;
        RECT  11.450 0.990 12.140 1.220 ;
        RECT  11.895 2.565 12.140 2.795 ;
        RECT  11.680 1.530 11.910 2.300 ;
        RECT  11.375 2.070 11.680 2.300 ;
        RECT  11.220 0.990 11.450 1.830 ;
        RECT  11.145 2.070 11.375 2.995 ;
        RECT  10.655 1.600 11.220 1.830 ;
        RECT  9.610 2.765 11.145 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.070 2.300 10.775 2.530 ;
        RECT  10.070 0.990 10.760 1.220 ;
        RECT  8.955 3.225 10.440 3.455 ;
        RECT  9.840 0.465 10.070 2.530 ;
        RECT  8.405 0.465 9.840 0.695 ;
        RECT  9.380 0.925 9.610 2.995 ;
        RECT  8.875 1.475 9.105 2.500 ;
        RECT  8.725 2.730 8.955 3.455 ;
        RECT  8.865 1.475 8.875 1.705 ;
        RECT  8.765 2.270 8.875 2.500 ;
        RECT  8.635 0.925 8.865 1.705 ;
        RECT  7.480 2.730 8.725 2.960 ;
        RECT  7.720 1.475 8.635 1.705 ;
        RECT  8.175 0.465 8.405 1.245 ;
        RECT  8.050 1.935 8.390 2.470 ;
        RECT  7.330 1.015 8.175 1.245 ;
        RECT  6.805 2.240 8.050 2.470 ;
        RECT  7.380 1.475 7.720 1.890 ;
        RECT  7.250 2.730 7.480 3.250 ;
        RECT  7.100 0.465 7.330 1.245 ;
        RECT  6.170 3.020 7.250 3.250 ;
        RECT  4.820 0.465 7.100 0.695 ;
        RECT  6.755 2.240 6.805 2.650 ;
        RECT  6.525 0.935 6.755 2.650 ;
        RECT  5.940 0.975 6.155 2.630 ;
        RECT  5.925 0.975 5.940 3.210 ;
        RECT  5.745 0.975 5.925 1.210 ;
        RECT  5.710 2.390 5.925 3.210 ;
        RECT  2.675 2.980 5.710 3.210 ;
        RECT  5.440 1.615 5.695 1.955 ;
        RECT  5.210 0.925 5.440 2.750 ;
        RECT  5.105 0.925 5.210 1.265 ;
        RECT  5.095 2.520 5.210 2.750 ;
        RECT  4.800 1.770 4.975 2.110 ;
        RECT  4.590 0.465 4.820 0.925 ;
        RECT  4.570 1.155 4.800 2.670 ;
        RECT  3.175 0.695 4.590 0.925 ;
        RECT  3.710 1.155 4.570 1.385 ;
        RECT  3.780 2.440 4.570 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.465 2.675 3.210 ;
        RECT  2.060 0.465 2.445 0.695 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFD0BWP7T

MACRO EDFD1BWP7T
    CLASS CORE ;
    FOREIGN EDFD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.0304 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.075 13.300 2.560 ;
        RECT  12.885 1.075 13.020 1.305 ;
        RECT  12.600 2.330 13.020 2.560 ;
        RECT  12.655 0.920 12.885 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.470 14.420 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.660 0.810 ;
        RECT  10.530 -0.235 13.320 0.235 ;
        RECT  10.300 -0.235 10.530 0.520 ;
        RECT  7.945 -0.235 10.300 0.235 ;
        RECT  7.715 -0.235 7.945 0.785 ;
        RECT  4.360 -0.235 7.715 0.235 ;
        RECT  4.020 -0.235 4.360 0.465 ;
        RECT  3.660 -0.235 4.020 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 3.685 14.560 4.155 ;
        RECT  13.320 3.250 13.660 4.155 ;
        RECT  11.515 3.685 13.320 4.155 ;
        RECT  11.170 3.225 11.515 4.155 ;
        RECT  8.185 3.685 11.170 4.155 ;
        RECT  7.825 3.190 8.185 4.155 ;
        RECT  4.680 3.685 7.825 4.155 ;
        RECT  4.340 3.455 4.680 4.155 ;
        RECT  3.620 3.685 4.340 4.155 ;
        RECT  3.280 3.455 3.620 4.155 ;
        RECT  1.250 3.685 3.280 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.020 ;
        RECT  12.370 2.790 13.615 3.020 ;
        RECT  10.990 0.465 12.580 0.695 ;
        RECT  12.180 1.020 12.370 3.020 ;
        RECT  12.140 1.020 12.180 3.380 ;
        RECT  11.450 1.020 12.140 1.250 ;
        RECT  11.950 2.565 12.140 3.380 ;
        RECT  11.680 1.530 11.910 2.300 ;
        RECT  11.375 2.070 11.680 2.300 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  11.145 2.070 11.375 2.995 ;
        RECT  10.655 1.600 11.220 1.830 ;
        RECT  9.610 2.765 11.145 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.070 2.300 10.775 2.530 ;
        RECT  10.070 0.990 10.760 1.220 ;
        RECT  8.955 3.225 10.440 3.455 ;
        RECT  9.840 0.465 10.070 2.530 ;
        RECT  8.405 0.465 9.840 0.695 ;
        RECT  9.380 0.925 9.610 2.995 ;
        RECT  8.875 1.475 9.105 2.500 ;
        RECT  8.725 2.730 8.955 3.455 ;
        RECT  8.865 1.475 8.875 1.705 ;
        RECT  8.765 2.270 8.875 2.500 ;
        RECT  8.635 0.925 8.865 1.705 ;
        RECT  7.480 2.730 8.725 2.960 ;
        RECT  7.720 1.475 8.635 1.705 ;
        RECT  8.175 0.465 8.405 1.245 ;
        RECT  8.050 1.935 8.390 2.470 ;
        RECT  7.330 1.015 8.175 1.245 ;
        RECT  6.805 2.240 8.050 2.470 ;
        RECT  7.380 1.475 7.720 1.890 ;
        RECT  7.250 2.730 7.480 3.250 ;
        RECT  7.100 0.465 7.330 1.245 ;
        RECT  6.170 3.020 7.250 3.250 ;
        RECT  4.820 0.465 7.100 0.695 ;
        RECT  6.755 2.240 6.805 2.650 ;
        RECT  6.525 0.935 6.755 2.650 ;
        RECT  5.940 0.975 6.155 2.630 ;
        RECT  5.925 0.975 5.940 3.210 ;
        RECT  5.745 0.975 5.925 1.210 ;
        RECT  5.710 2.390 5.925 3.210 ;
        RECT  2.675 2.980 5.710 3.210 ;
        RECT  5.440 1.615 5.695 1.955 ;
        RECT  5.210 0.925 5.440 2.750 ;
        RECT  5.105 0.925 5.210 1.265 ;
        RECT  5.095 2.520 5.210 2.750 ;
        RECT  4.800 1.770 4.975 2.110 ;
        RECT  4.590 0.465 4.820 0.925 ;
        RECT  4.570 1.155 4.800 2.670 ;
        RECT  3.175 0.695 4.590 0.925 ;
        RECT  3.710 1.155 4.570 1.385 ;
        RECT  3.780 2.440 4.570 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.465 2.675 3.210 ;
        RECT  2.060 0.465 2.445 0.695 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFD1BWP7T

MACRO EDFD2BWP7T
    CLASS CORE ;
    FOREIGN EDFD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.860 2.330 13.900 2.560 ;
        RECT  13.580 0.465 13.860 2.560 ;
        RECT  13.560 2.330 13.580 2.560 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.035 15.540 2.615 ;
        RECT  15.260 0.465 15.285 3.310 ;
        RECT  15.055 0.465 15.260 1.315 ;
        RECT  15.055 2.360 15.260 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.340 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.315 ;
        RECT  14.565 -0.235 15.775 0.235 ;
        RECT  14.335 -0.235 14.565 1.290 ;
        RECT  13.125 -0.235 14.335 0.235 ;
        RECT  12.895 -0.235 13.125 0.925 ;
        RECT  11.405 -0.235 12.895 0.235 ;
        RECT  11.175 -0.235 11.405 0.520 ;
        RECT  7.945 -0.235 11.175 0.235 ;
        RECT  7.715 -0.235 7.945 0.785 ;
        RECT  4.360 -0.235 7.715 0.235 ;
        RECT  4.020 -0.235 4.360 0.465 ;
        RECT  3.660 -0.235 4.020 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.250 -0.235 3.320 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.245 16.005 4.155 ;
        RECT  14.620 3.685 15.775 4.155 ;
        RECT  14.280 3.250 14.620 4.155 ;
        RECT  12.975 3.685 14.280 4.155 ;
        RECT  12.635 3.250 12.975 4.155 ;
        RECT  11.515 3.685 12.635 4.155 ;
        RECT  11.170 3.225 11.515 4.155 ;
        RECT  8.185 3.685 11.170 4.155 ;
        RECT  7.825 3.190 8.185 4.155 ;
        RECT  4.680 3.685 7.825 4.155 ;
        RECT  4.340 3.455 4.680 4.155 ;
        RECT  3.620 3.685 4.340 4.155 ;
        RECT  3.280 3.455 3.620 4.155 ;
        RECT  1.250 3.685 3.280 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.580 1.600 14.810 3.020 ;
        RECT  13.145 2.790 14.580 3.020 ;
        RECT  12.915 1.265 13.145 3.020 ;
        RECT  12.325 1.265 12.915 1.495 ;
        RECT  12.180 2.565 12.915 2.795 ;
        RECT  11.865 0.500 12.660 0.730 ;
        RECT  12.095 0.965 12.325 1.495 ;
        RECT  11.950 2.565 12.180 3.380 ;
        RECT  10.940 1.265 12.095 1.495 ;
        RECT  11.595 1.780 12.020 2.010 ;
        RECT  11.635 0.500 11.865 1.035 ;
        RECT  10.280 0.805 11.635 1.035 ;
        RECT  11.365 1.780 11.595 2.995 ;
        RECT  9.610 2.765 11.365 2.995 ;
        RECT  10.710 1.265 10.940 1.900 ;
        RECT  10.280 2.300 10.775 2.530 ;
        RECT  8.955 3.225 10.440 3.455 ;
        RECT  10.050 0.465 10.280 2.530 ;
        RECT  8.405 0.465 10.050 0.695 ;
        RECT  9.380 0.925 9.610 2.995 ;
        RECT  8.875 1.475 9.105 2.500 ;
        RECT  8.725 2.730 8.955 3.455 ;
        RECT  8.865 1.475 8.875 1.705 ;
        RECT  8.765 2.270 8.875 2.500 ;
        RECT  8.635 0.925 8.865 1.705 ;
        RECT  7.480 2.730 8.725 2.960 ;
        RECT  7.720 1.475 8.635 1.705 ;
        RECT  8.175 0.465 8.405 1.245 ;
        RECT  8.050 1.935 8.390 2.470 ;
        RECT  7.330 1.015 8.175 1.245 ;
        RECT  6.805 2.240 8.050 2.470 ;
        RECT  7.380 1.475 7.720 1.890 ;
        RECT  7.250 2.730 7.480 3.250 ;
        RECT  7.100 0.465 7.330 1.245 ;
        RECT  6.170 3.020 7.250 3.250 ;
        RECT  4.820 0.465 7.100 0.695 ;
        RECT  6.755 2.240 6.805 2.650 ;
        RECT  6.525 0.935 6.755 2.650 ;
        RECT  5.940 0.975 6.155 2.630 ;
        RECT  5.925 0.975 5.940 3.210 ;
        RECT  5.745 0.975 5.925 1.210 ;
        RECT  5.710 2.390 5.925 3.210 ;
        RECT  2.675 2.980 5.710 3.210 ;
        RECT  5.440 1.615 5.695 1.955 ;
        RECT  5.210 0.925 5.440 2.750 ;
        RECT  5.105 0.925 5.210 1.265 ;
        RECT  5.095 2.520 5.210 2.750 ;
        RECT  4.800 1.770 4.975 2.110 ;
        RECT  4.590 0.465 4.820 0.925 ;
        RECT  4.570 1.155 4.800 2.670 ;
        RECT  3.175 0.695 4.590 0.925 ;
        RECT  3.710 1.155 4.570 1.385 ;
        RECT  3.780 2.440 4.570 2.670 ;
        RECT  2.945 0.695 3.175 2.270 ;
        RECT  2.445 0.465 2.675 3.210 ;
        RECT  2.060 0.465 2.445 0.695 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFD2BWP7T

MACRO EDFKCND0BWP7T
    CLASS CORE ;
    FOREIGN EDFKCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 0.5938 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.215 0.950 15.540 2.710 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.140 0.965 14.420 2.560 ;
        RECT  13.845 0.965 14.140 1.305 ;
        RECT  13.720 2.330 14.140 2.560 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.610 0.705 1.845 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2322 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 2.000 2.450 2.230 ;
        RECT  1.820 1.765 2.100 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.125 2.330 6.580 2.710 ;
        RECT  5.895 1.765 6.125 2.710 ;
        RECT  5.740 1.765 5.895 2.150 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.210 4.420 2.210 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.445 -0.235 15.680 0.235 ;
        RECT  15.215 -0.235 15.445 0.545 ;
        RECT  9.495 -0.235 15.215 0.235 ;
        RECT  9.265 -0.235 9.495 0.520 ;
        RECT  6.180 -0.235 9.265 0.235 ;
        RECT  5.840 -0.235 6.180 0.465 ;
        RECT  5.105 -0.235 5.840 0.235 ;
        RECT  4.760 -0.235 5.105 0.465 ;
        RECT  0.475 -0.235 4.760 0.235 ;
        RECT  0.230 -0.235 0.475 0.930 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.780 3.685 15.680 4.155 ;
        RECT  14.440 3.290 14.780 4.155 ;
        RECT  13.445 3.685 14.440 4.155 ;
        RECT  13.100 3.455 13.445 4.155 ;
        RECT  9.720 3.685 13.100 4.155 ;
        RECT  9.360 3.190 9.720 4.155 ;
        RECT  6.285 3.685 9.360 4.155 ;
        RECT  5.945 3.455 6.285 4.155 ;
        RECT  4.230 3.685 5.945 4.155 ;
        RECT  3.885 3.455 4.230 4.155 ;
        RECT  1.195 3.685 3.885 4.155 ;
        RECT  0.945 2.855 1.195 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.755 0.465 14.985 3.020 ;
        RECT  12.055 0.465 14.755 0.695 ;
        RECT  14.095 2.790 14.755 3.020 ;
        RECT  13.850 2.790 14.095 3.220 ;
        RECT  13.490 1.580 13.900 1.970 ;
        RECT  12.835 2.990 13.850 3.220 ;
        RECT  13.260 0.965 13.490 2.760 ;
        RECT  12.570 0.965 13.260 1.195 ;
        RECT  13.000 2.530 13.260 2.760 ;
        RECT  12.800 1.530 13.030 2.300 ;
        RECT  12.605 2.990 12.835 3.455 ;
        RECT  12.355 2.070 12.800 2.300 ;
        RECT  10.380 3.225 12.605 3.455 ;
        RECT  12.340 0.965 12.570 1.830 ;
        RECT  12.125 2.070 12.355 2.995 ;
        RECT  12.010 1.600 12.340 1.830 ;
        RECT  11.135 2.765 12.125 2.995 ;
        RECT  11.825 0.465 12.055 1.275 ;
        RECT  11.595 2.305 11.845 2.535 ;
        RECT  11.365 0.465 11.595 2.535 ;
        RECT  9.955 0.465 11.365 0.695 ;
        RECT  10.905 0.925 11.135 2.995 ;
        RECT  10.415 1.290 10.535 2.500 ;
        RECT  10.305 0.935 10.415 2.500 ;
        RECT  10.150 2.730 10.380 3.455 ;
        RECT  10.185 0.935 10.305 1.520 ;
        RECT  10.130 2.270 10.305 2.500 ;
        RECT  9.345 1.290 10.185 1.520 ;
        RECT  9.025 2.730 10.150 2.960 ;
        RECT  9.890 1.750 10.075 1.980 ;
        RECT  9.725 0.465 9.955 1.060 ;
        RECT  9.660 1.750 9.890 2.475 ;
        RECT  8.895 0.830 9.725 1.060 ;
        RECT  8.465 2.245 9.660 2.475 ;
        RECT  9.115 1.290 9.345 1.965 ;
        RECT  8.790 2.730 9.025 3.425 ;
        RECT  8.665 0.465 8.895 1.060 ;
        RECT  7.175 3.195 8.790 3.425 ;
        RECT  8.510 0.465 8.665 0.695 ;
        RECT  8.435 2.245 8.465 2.845 ;
        RECT  8.205 0.935 8.435 2.845 ;
        RECT  7.745 0.500 7.975 2.790 ;
        RECT  6.655 0.500 7.745 0.730 ;
        RECT  7.515 2.450 7.745 2.790 ;
        RECT  7.285 1.615 7.515 1.955 ;
        RECT  7.055 1.085 7.285 2.765 ;
        RECT  6.935 2.995 7.175 3.425 ;
        RECT  6.830 1.085 7.055 1.440 ;
        RECT  6.815 2.425 7.055 2.765 ;
        RECT  3.565 2.995 6.935 3.225 ;
        RECT  6.585 1.750 6.805 2.090 ;
        RECT  6.425 0.500 6.655 0.925 ;
        RECT  6.355 1.155 6.585 2.090 ;
        RECT  4.965 0.695 6.425 0.925 ;
        RECT  5.510 1.155 6.355 1.385 ;
        RECT  5.510 2.410 5.665 2.765 ;
        RECT  5.280 1.155 5.510 2.765 ;
        RECT  4.735 0.695 4.965 2.765 ;
        RECT  3.615 0.695 4.735 0.925 ;
        RECT  3.385 0.695 3.615 2.750 ;
        RECT  3.335 2.995 3.565 3.335 ;
        RECT  2.550 0.775 3.385 1.005 ;
        RECT  2.350 2.520 3.385 2.750 ;
        RECT  2.835 1.235 3.065 1.730 ;
        RECT  1.575 1.235 2.835 1.465 ;
        RECT  1.335 1.235 1.575 2.625 ;
        RECT  1.195 1.235 1.335 1.465 ;
        RECT  0.470 2.385 1.335 2.625 ;
        RECT  0.950 0.610 1.195 1.465 ;
        RECT  0.230 2.385 0.470 3.165 ;
    END
END EDFKCND0BWP7T

MACRO EDFKCND1BWP7T
    CLASS CORE ;
    FOREIGN EDFKCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.3926 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.510 2.380 6.070 2.740 ;
        RECT  5.510 0.925 5.545 1.610 ;
        RECT  5.315 0.925 5.510 2.740 ;
        RECT  5.280 1.395 5.315 2.740 ;
        RECT  5.030 2.380 5.280 2.740 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.215 0.465 15.540 3.345 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.610 0.705 1.845 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2322 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 2.000 2.305 2.230 ;
        RECT  1.820 1.765 2.100 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.770 6.590 2.150 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.160 4.340 2.210 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.215 -0.235 15.680 0.235 ;
        RECT  12.985 -0.235 13.215 0.575 ;
        RECT  9.915 -0.235 12.985 0.235 ;
        RECT  9.685 -0.235 9.915 0.520 ;
        RECT  6.585 -0.235 9.685 0.235 ;
        RECT  6.245 -0.235 6.585 0.465 ;
        RECT  4.625 -0.235 6.245 0.235 ;
        RECT  4.395 -0.235 4.625 0.750 ;
        RECT  0.475 -0.235 4.395 0.235 ;
        RECT  0.230 -0.235 0.475 0.945 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.720 3.685 15.680 4.155 ;
        RECT  14.375 3.455 14.720 4.155 ;
        RECT  13.410 3.685 14.375 4.155 ;
        RECT  13.070 3.455 13.410 4.155 ;
        RECT  10.405 3.685 13.070 4.155 ;
        RECT  10.045 3.190 10.405 4.155 ;
        RECT  7.090 3.685 10.045 4.155 ;
        RECT  6.750 3.455 7.090 4.155 ;
        RECT  6.075 3.685 6.750 4.155 ;
        RECT  5.735 3.455 6.075 4.155 ;
        RECT  3.800 3.685 5.735 4.155 ;
        RECT  3.455 3.455 3.800 4.155 ;
        RECT  1.195 3.685 3.455 4.155 ;
        RECT  0.945 2.855 1.195 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.755 0.490 14.985 2.990 ;
        RECT  13.675 0.490 14.755 0.720 ;
        RECT  12.870 2.760 14.755 2.990 ;
        RECT  14.295 1.265 14.525 2.530 ;
        RECT  14.135 1.265 14.295 1.495 ;
        RECT  13.830 2.300 14.295 2.530 ;
        RECT  13.905 0.960 14.135 1.495 ;
        RECT  12.990 1.265 13.905 1.495 ;
        RECT  13.475 1.775 13.790 2.015 ;
        RECT  13.445 0.490 13.675 1.035 ;
        RECT  13.245 1.775 13.475 2.300 ;
        RECT  12.535 0.805 13.445 1.035 ;
        RECT  12.075 2.060 13.245 2.300 ;
        RECT  12.650 1.265 12.990 1.830 ;
        RECT  12.510 2.705 12.870 2.990 ;
        RECT  12.305 0.465 12.535 1.035 ;
        RECT  11.615 3.225 12.320 3.455 ;
        RECT  10.375 0.465 12.305 0.695 ;
        RECT  11.845 0.925 12.075 2.990 ;
        RECT  11.325 0.925 11.845 1.155 ;
        RECT  11.385 1.390 11.615 3.455 ;
        RECT  11.265 1.390 11.385 1.730 ;
        RECT  9.765 2.730 11.385 2.960 ;
        RECT  11.035 2.265 11.155 2.500 ;
        RECT  10.945 1.215 11.035 2.500 ;
        RECT  10.805 0.925 10.945 2.500 ;
        RECT  10.605 0.925 10.805 1.445 ;
        RECT  9.905 1.215 10.605 1.445 ;
        RECT  10.495 1.695 10.575 2.035 ;
        RECT  10.265 1.695 10.495 2.290 ;
        RECT  10.145 0.465 10.375 0.985 ;
        RECT  9.150 2.060 10.265 2.290 ;
        RECT  9.455 0.755 10.145 0.985 ;
        RECT  9.675 1.215 9.905 1.815 ;
        RECT  9.535 2.730 9.765 3.250 ;
        RECT  8.625 3.020 9.535 3.250 ;
        RECT  9.225 0.465 9.455 0.985 ;
        RECT  7.045 0.465 9.225 0.695 ;
        RECT  8.995 2.060 9.150 2.785 ;
        RECT  8.765 0.935 8.995 2.785 ;
        RECT  8.395 0.925 8.500 2.730 ;
        RECT  8.270 0.925 8.395 3.455 ;
        RECT  8.045 0.925 8.270 1.265 ;
        RECT  8.165 2.500 8.270 3.455 ;
        RECT  8.155 2.995 8.165 3.455 ;
        RECT  4.575 2.995 8.155 3.225 ;
        RECT  7.850 1.585 8.040 1.925 ;
        RECT  7.795 1.585 7.850 2.740 ;
        RECT  7.565 0.940 7.795 2.740 ;
        RECT  7.290 0.940 7.565 1.170 ;
        RECT  7.050 1.490 7.335 1.830 ;
        RECT  6.820 1.155 7.050 2.740 ;
        RECT  6.815 0.465 7.045 0.925 ;
        RECT  5.950 1.155 6.820 1.385 ;
        RECT  6.300 2.400 6.820 2.740 ;
        RECT  6.005 0.695 6.815 0.925 ;
        RECT  5.775 0.465 6.005 0.925 ;
        RECT  5.085 0.465 5.775 0.695 ;
        RECT  5.010 0.465 5.085 1.240 ;
        RECT  4.855 0.465 5.010 1.930 ;
        RECT  4.800 1.030 4.855 1.930 ;
        RECT  4.780 1.030 4.800 2.670 ;
        RECT  4.570 1.590 4.780 2.670 ;
        RECT  4.235 2.995 4.575 3.455 ;
        RECT  3.155 2.440 4.570 2.670 ;
        RECT  2.835 2.995 4.235 3.225 ;
        RECT  3.295 0.775 3.525 2.190 ;
        RECT  2.550 0.775 3.295 1.005 ;
        RECT  2.800 1.960 3.295 2.190 ;
        RECT  2.835 1.235 3.065 1.730 ;
        RECT  1.575 1.235 2.835 1.465 ;
        RECT  2.800 2.995 2.835 3.355 ;
        RECT  2.570 1.960 2.800 3.355 ;
        RECT  2.300 3.010 2.570 3.355 ;
        RECT  1.335 1.235 1.575 2.625 ;
        RECT  1.195 1.235 1.335 1.465 ;
        RECT  0.470 2.385 1.335 2.625 ;
        RECT  0.950 0.625 1.195 1.465 ;
        RECT  0.230 2.385 0.470 3.165 ;
    END
END EDFKCND1BWP7T

MACRO EDFKCND2BWP7T
    CLASS CORE ;
    FOREIGN EDFKCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.405 1.050 16.660 2.625 ;
        RECT  16.380 0.465 16.405 3.310 ;
        RECT  16.175 0.465 16.380 1.290 ;
        RECT  16.175 2.350 16.380 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.980 2.300 15.020 2.530 ;
        RECT  14.680 0.465 14.980 2.530 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.610 0.705 1.845 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2322 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 2.000 2.450 2.230 ;
        RECT  1.820 1.765 2.100 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.770 6.020 2.150 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.160 4.340 2.210 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.125 -0.235 17.360 0.235 ;
        RECT  16.895 -0.235 17.125 1.290 ;
        RECT  15.685 -0.235 16.895 0.235 ;
        RECT  15.455 -0.235 15.685 1.215 ;
        RECT  12.775 -0.235 15.455 0.235 ;
        RECT  12.545 -0.235 12.775 0.520 ;
        RECT  9.355 -0.235 12.545 0.235 ;
        RECT  9.125 -0.235 9.355 0.520 ;
        RECT  6.020 -0.235 9.125 0.235 ;
        RECT  5.680 -0.235 6.020 0.465 ;
        RECT  5.105 -0.235 5.680 0.235 ;
        RECT  4.760 -0.235 5.105 0.465 ;
        RECT  0.475 -0.235 4.760 0.235 ;
        RECT  0.230 -0.235 0.475 0.955 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.125 3.685 17.360 4.155 ;
        RECT  16.895 2.245 17.125 4.155 ;
        RECT  15.740 3.685 16.895 4.155 ;
        RECT  15.400 3.250 15.740 4.155 ;
        RECT  14.240 3.685 15.400 4.155 ;
        RECT  13.895 3.455 14.240 4.155 ;
        RECT  12.930 3.685 13.895 4.155 ;
        RECT  12.590 3.455 12.930 4.155 ;
        RECT  9.720 3.685 12.590 4.155 ;
        RECT  9.360 3.190 9.720 4.155 ;
        RECT  6.285 3.685 9.360 4.155 ;
        RECT  5.945 3.455 6.285 4.155 ;
        RECT  4.230 3.685 5.945 4.155 ;
        RECT  3.885 3.455 4.230 4.155 ;
        RECT  1.195 3.685 3.885 4.155 ;
        RECT  0.945 2.855 1.195 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.695 1.655 16.120 1.885 ;
        RECT  15.465 1.655 15.695 2.990 ;
        RECT  14.360 2.760 15.465 2.990 ;
        RECT  14.130 0.490 14.360 2.990 ;
        RECT  13.235 0.490 14.130 0.720 ;
        RECT  12.270 2.760 14.130 2.990 ;
        RECT  13.695 1.265 13.900 2.530 ;
        RECT  13.670 0.960 13.695 2.530 ;
        RECT  13.465 0.960 13.670 1.535 ;
        RECT  13.385 2.300 13.670 2.530 ;
        RECT  12.470 1.305 13.465 1.535 ;
        RECT  13.005 0.490 13.235 1.075 ;
        RECT  13.100 1.780 13.210 2.010 ;
        RECT  12.870 1.780 13.100 2.300 ;
        RECT  11.960 0.845 13.005 1.075 ;
        RECT  11.475 2.070 12.870 2.300 ;
        RECT  12.130 1.305 12.470 1.830 ;
        RECT  11.910 2.705 12.270 2.990 ;
        RECT  11.730 0.465 11.960 1.075 ;
        RECT  10.935 3.225 11.890 3.455 ;
        RECT  9.815 0.465 11.730 0.695 ;
        RECT  11.455 2.070 11.475 2.990 ;
        RECT  11.225 0.925 11.455 2.990 ;
        RECT  10.890 0.925 11.225 1.155 ;
        RECT  10.705 1.390 10.935 3.455 ;
        RECT  8.960 2.730 10.705 2.960 ;
        RECT  10.275 1.215 10.475 2.500 ;
        RECT  10.245 0.935 10.275 2.500 ;
        RECT  10.045 0.935 10.245 1.445 ;
        RECT  10.130 2.270 10.245 2.500 ;
        RECT  9.345 1.215 10.045 1.445 ;
        RECT  9.805 1.695 10.015 2.035 ;
        RECT  9.585 0.465 9.815 0.985 ;
        RECT  9.575 1.695 9.805 2.500 ;
        RECT  8.895 0.755 9.585 0.985 ;
        RECT  8.465 2.270 9.575 2.500 ;
        RECT  9.115 1.215 9.345 2.020 ;
        RECT  8.730 2.730 8.960 3.250 ;
        RECT  8.665 0.465 8.895 0.985 ;
        RECT  7.940 3.020 8.730 3.250 ;
        RECT  6.490 0.465 8.665 0.695 ;
        RECT  8.435 2.270 8.465 2.785 ;
        RECT  8.205 0.935 8.435 2.785 ;
        RECT  7.745 0.980 7.975 2.730 ;
        RECT  7.430 0.980 7.745 1.210 ;
        RECT  7.590 2.500 7.745 2.730 ;
        RECT  7.360 2.500 7.590 3.225 ;
        RECT  7.130 1.585 7.515 1.925 ;
        RECT  3.065 2.995 7.360 3.225 ;
        RECT  6.900 0.925 7.130 2.765 ;
        RECT  6.730 0.925 6.900 1.155 ;
        RECT  6.815 2.425 6.900 2.765 ;
        RECT  6.480 1.750 6.670 2.090 ;
        RECT  6.260 0.465 6.490 0.925 ;
        RECT  6.250 1.155 6.480 2.740 ;
        RECT  4.845 0.695 6.260 0.925 ;
        RECT  5.280 1.155 6.250 1.385 ;
        RECT  5.440 2.510 6.250 2.740 ;
        RECT  4.615 0.695 4.845 2.670 ;
        RECT  3.555 2.440 4.615 2.670 ;
        RECT  3.385 0.775 3.615 2.190 ;
        RECT  2.550 0.775 3.385 1.005 ;
        RECT  3.065 1.960 3.385 2.190 ;
        RECT  2.835 1.235 3.065 1.730 ;
        RECT  2.835 1.960 3.065 3.225 ;
        RECT  1.575 1.235 2.835 1.465 ;
        RECT  2.405 2.760 2.835 3.105 ;
        RECT  1.335 1.235 1.575 2.625 ;
        RECT  1.195 1.235 1.335 1.465 ;
        RECT  0.470 2.385 1.335 2.625 ;
        RECT  0.950 0.660 1.195 1.465 ;
        RECT  0.230 2.385 0.470 3.165 ;
    END
END EDFKCND2BWP7T

MACRO EDFKCNQD1BWP7T
    CLASS CORE ;
    FOREIGN EDFKCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.120 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.655 0.470 14.980 3.265 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.610 0.705 1.845 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2322 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 2.000 2.450 2.230 ;
        RECT  1.820 1.765 2.100 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.770 6.020 2.150 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.160 4.340 2.210 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.705 -0.235 15.120 0.235 ;
        RECT  12.475 -0.235 12.705 0.520 ;
        RECT  9.285 -0.235 12.475 0.235 ;
        RECT  9.055 -0.235 9.285 0.520 ;
        RECT  5.850 -0.235 9.055 0.235 ;
        RECT  5.510 -0.235 5.850 0.465 ;
        RECT  4.850 -0.235 5.510 0.235 ;
        RECT  4.505 -0.235 4.850 0.465 ;
        RECT  0.475 -0.235 4.505 0.235 ;
        RECT  0.230 -0.235 0.475 0.950 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.180 3.685 15.120 4.155 ;
        RECT  13.835 3.455 14.180 4.155 ;
        RECT  12.860 3.685 13.835 4.155 ;
        RECT  12.520 3.455 12.860 4.155 ;
        RECT  9.650 3.685 12.520 4.155 ;
        RECT  9.290 3.190 9.650 4.155 ;
        RECT  6.270 3.685 9.290 4.155 ;
        RECT  5.930 3.455 6.270 4.155 ;
        RECT  4.185 3.685 5.930 4.155 ;
        RECT  3.840 3.455 4.185 4.155 ;
        RECT  1.195 3.685 3.840 4.155 ;
        RECT  0.945 2.855 1.195 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.090 0.465 14.320 2.990 ;
        RECT  13.165 0.465 14.090 0.695 ;
        RECT  12.200 2.760 14.090 2.990 ;
        RECT  13.625 1.265 13.830 2.530 ;
        RECT  13.600 0.960 13.625 2.530 ;
        RECT  13.395 0.960 13.600 1.495 ;
        RECT  13.315 2.300 13.600 2.530 ;
        RECT  12.400 1.265 13.395 1.495 ;
        RECT  12.935 0.465 13.165 1.035 ;
        RECT  12.855 1.725 13.085 2.300 ;
        RECT  11.890 0.805 12.935 1.035 ;
        RECT  11.405 2.070 12.855 2.300 ;
        RECT  12.060 1.265 12.400 1.830 ;
        RECT  11.840 2.705 12.200 2.990 ;
        RECT  11.660 0.465 11.890 1.035 ;
        RECT  10.865 3.225 11.820 3.455 ;
        RECT  9.745 0.465 11.660 0.695 ;
        RECT  11.385 2.070 11.405 2.990 ;
        RECT  11.155 0.925 11.385 2.990 ;
        RECT  10.820 0.925 11.155 1.155 ;
        RECT  10.635 1.390 10.865 3.455 ;
        RECT  8.890 2.730 10.635 2.960 ;
        RECT  10.205 1.215 10.405 2.500 ;
        RECT  10.175 0.935 10.205 2.500 ;
        RECT  9.975 0.935 10.175 1.445 ;
        RECT  10.060 2.270 10.175 2.500 ;
        RECT  9.275 1.215 9.975 1.445 ;
        RECT  9.735 1.695 9.945 2.035 ;
        RECT  9.515 0.465 9.745 0.985 ;
        RECT  9.505 1.695 9.735 2.500 ;
        RECT  8.825 0.755 9.515 0.985 ;
        RECT  8.395 2.270 9.505 2.500 ;
        RECT  9.045 1.215 9.275 2.020 ;
        RECT  8.660 2.730 8.890 3.250 ;
        RECT  8.595 0.465 8.825 0.985 ;
        RECT  7.870 3.020 8.660 3.250 ;
        RECT  6.310 0.465 8.595 0.695 ;
        RECT  8.365 2.270 8.395 2.785 ;
        RECT  8.135 0.935 8.365 2.785 ;
        RECT  7.675 0.980 7.905 2.615 ;
        RECT  7.360 0.980 7.675 1.210 ;
        RECT  7.520 2.385 7.675 2.615 ;
        RECT  7.290 2.385 7.520 3.225 ;
        RECT  7.060 1.585 7.445 1.925 ;
        RECT  4.975 2.995 7.290 3.225 ;
        RECT  6.830 0.925 7.060 2.765 ;
        RECT  6.715 0.925 6.830 1.265 ;
        RECT  6.745 2.425 6.830 2.765 ;
        RECT  6.480 1.750 6.600 2.090 ;
        RECT  6.250 1.155 6.480 2.740 ;
        RECT  6.080 0.465 6.310 0.925 ;
        RECT  5.075 1.155 6.250 1.385 ;
        RECT  5.175 2.510 6.250 2.740 ;
        RECT  4.845 0.695 6.080 0.925 ;
        RECT  4.635 2.995 4.975 3.455 ;
        RECT  4.615 0.695 4.845 2.670 ;
        RECT  3.065 2.995 4.635 3.225 ;
        RECT  3.555 2.440 4.615 2.670 ;
        RECT  3.385 0.775 3.615 2.190 ;
        RECT  2.550 0.775 3.385 1.005 ;
        RECT  3.065 1.960 3.385 2.190 ;
        RECT  2.835 1.235 3.065 1.730 ;
        RECT  2.835 1.960 3.065 3.225 ;
        RECT  1.575 1.235 2.835 1.465 ;
        RECT  2.500 2.955 2.835 3.225 ;
        RECT  1.335 1.235 1.575 2.625 ;
        RECT  1.195 1.235 1.335 1.465 ;
        RECT  0.470 2.385 1.335 2.625 ;
        RECT  0.950 0.660 1.195 1.465 ;
        RECT  0.230 2.385 0.470 3.165 ;
    END
END EDFKCNQD1BWP7T

MACRO EDFKCNQD2BWP7T
    CLASS CORE ;
    FOREIGN EDFKCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.070 15.540 2.730 ;
        RECT  15.260 0.465 15.285 3.385 ;
        RECT  15.055 0.465 15.260 1.305 ;
        RECT  15.055 2.370 15.260 3.385 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.610 0.705 1.845 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2322 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 2.000 2.450 2.230 ;
        RECT  1.820 1.765 2.100 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.125 2.330 6.580 2.710 ;
        RECT  5.895 1.765 6.125 2.710 ;
        RECT  5.740 1.765 5.895 2.150 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.210 4.420 2.210 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.300 ;
        RECT  14.525 -0.235 15.775 0.235 ;
        RECT  14.295 -0.235 14.525 0.630 ;
        RECT  12.660 -0.235 14.295 0.235 ;
        RECT  12.430 -0.235 12.660 0.535 ;
        RECT  9.600 -0.235 12.430 0.235 ;
        RECT  9.260 -0.235 9.600 0.465 ;
        RECT  6.060 -0.235 9.260 0.235 ;
        RECT  5.720 -0.235 6.060 0.465 ;
        RECT  5.105 -0.235 5.720 0.235 ;
        RECT  4.760 -0.235 5.105 0.465 ;
        RECT  0.475 -0.235 4.760 0.235 ;
        RECT  0.230 -0.235 0.475 0.930 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.245 16.005 4.155 ;
        RECT  14.580 3.685 15.775 4.155 ;
        RECT  14.235 3.455 14.580 4.155 ;
        RECT  13.185 3.685 14.235 4.155 ;
        RECT  12.955 3.400 13.185 4.155 ;
        RECT  9.830 3.685 12.955 4.155 ;
        RECT  9.470 3.190 9.830 4.155 ;
        RECT  6.285 3.685 9.470 4.155 ;
        RECT  5.945 3.455 6.285 4.155 ;
        RECT  4.230 3.685 5.945 4.155 ;
        RECT  3.885 3.455 4.230 4.155 ;
        RECT  1.195 3.685 3.885 4.155 ;
        RECT  0.945 2.855 1.195 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.595 0.860 14.825 3.125 ;
        RECT  14.065 0.860 14.595 1.090 ;
        RECT  12.725 2.895 14.595 3.125 ;
        RECT  14.110 1.320 14.340 2.600 ;
        RECT  13.605 1.320 14.110 1.550 ;
        RECT  13.740 2.370 14.110 2.600 ;
        RECT  13.835 0.505 14.065 1.090 ;
        RECT  13.145 0.505 13.835 0.735 ;
        RECT  13.375 0.965 13.605 1.550 ;
        RECT  13.130 1.780 13.470 2.300 ;
        RECT  12.820 1.320 13.375 1.550 ;
        RECT  12.915 0.505 13.145 1.090 ;
        RECT  12.265 2.070 13.130 2.300 ;
        RECT  12.165 0.860 12.915 1.090 ;
        RECT  12.590 1.320 12.820 1.830 ;
        RECT  12.495 2.895 12.725 3.455 ;
        RECT  12.120 1.600 12.590 1.830 ;
        RECT  10.490 3.225 12.495 3.455 ;
        RECT  12.035 2.070 12.265 2.995 ;
        RECT  11.935 0.860 12.165 1.275 ;
        RECT  11.245 2.765 12.035 2.995 ;
        RECT  11.705 2.195 11.805 2.535 ;
        RECT  11.475 0.465 11.705 2.535 ;
        RECT  10.065 0.465 11.475 0.695 ;
        RECT  11.015 0.925 11.245 2.995 ;
        RECT  10.525 1.290 10.645 2.500 ;
        RECT  10.415 0.935 10.525 2.500 ;
        RECT  10.260 2.730 10.490 3.455 ;
        RECT  10.295 0.935 10.415 1.520 ;
        RECT  10.240 2.270 10.415 2.500 ;
        RECT  9.455 1.290 10.295 1.520 ;
        RECT  9.105 2.730 10.260 2.960 ;
        RECT  10.000 1.750 10.185 1.980 ;
        RECT  9.835 0.465 10.065 1.060 ;
        RECT  9.770 1.750 10.000 2.475 ;
        RECT  8.975 0.830 9.835 1.060 ;
        RECT  8.545 2.245 9.770 2.475 ;
        RECT  9.225 1.290 9.455 1.965 ;
        RECT  8.870 2.730 9.105 3.425 ;
        RECT  8.745 0.465 8.975 1.060 ;
        RECT  7.175 3.195 8.870 3.425 ;
        RECT  8.590 0.465 8.745 0.695 ;
        RECT  8.515 2.245 8.545 2.845 ;
        RECT  8.285 0.935 8.515 2.845 ;
        RECT  7.825 0.465 8.055 2.880 ;
        RECT  7.510 0.465 7.825 0.730 ;
        RECT  7.595 2.470 7.825 2.880 ;
        RECT  7.285 1.615 7.515 1.955 ;
        RECT  6.545 0.465 7.510 0.695 ;
        RECT  7.055 0.925 7.285 2.765 ;
        RECT  6.935 2.995 7.175 3.425 ;
        RECT  6.830 0.925 7.055 1.265 ;
        RECT  6.815 2.425 7.055 2.765 ;
        RECT  3.765 2.995 6.935 3.225 ;
        RECT  6.585 1.750 6.805 2.090 ;
        RECT  6.355 1.155 6.585 2.090 ;
        RECT  6.315 0.465 6.545 0.925 ;
        RECT  5.510 1.155 6.355 1.385 ;
        RECT  4.965 0.695 6.315 0.925 ;
        RECT  5.510 2.410 5.665 2.765 ;
        RECT  5.280 1.155 5.510 2.765 ;
        RECT  4.735 0.695 4.965 2.720 ;
        RECT  3.615 0.695 4.735 0.925 ;
        RECT  3.420 2.440 3.765 3.225 ;
        RECT  3.385 0.695 3.615 2.190 ;
        RECT  2.550 0.775 3.385 1.005 ;
        RECT  2.980 1.960 3.385 2.190 ;
        RECT  2.835 1.235 3.065 1.730 ;
        RECT  2.750 1.960 2.980 3.270 ;
        RECT  1.575 1.235 2.835 1.465 ;
        RECT  2.490 2.925 2.750 3.270 ;
        RECT  1.335 1.235 1.575 2.625 ;
        RECT  1.195 1.235 1.335 1.465 ;
        RECT  0.470 2.385 1.335 2.625 ;
        RECT  0.950 0.610 1.195 1.465 ;
        RECT  0.230 2.385 0.470 3.165 ;
    END
END EDFKCNQD2BWP7T

MACRO EDFQD0BWP7T
    CLASS CORE ;
    FOREIGN EDFQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.530 0.555 13.860 3.085 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.345 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.045 -0.235 14.000 0.235 ;
        RECT  12.815 -0.235 13.045 0.865 ;
        RECT  11.495 -0.235 12.815 0.235 ;
        RECT  11.265 -0.235 11.495 0.665 ;
        RECT  8.110 -0.235 11.265 0.235 ;
        RECT  7.880 -0.235 8.110 0.785 ;
        RECT  4.415 -0.235 7.880 0.235 ;
        RECT  4.075 -0.235 4.415 0.465 ;
        RECT  3.715 -0.235 4.075 0.235 ;
        RECT  3.375 -0.235 3.715 0.465 ;
        RECT  1.250 -0.235 3.375 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.055 3.685 14.000 4.155 ;
        RECT  12.810 2.730 13.055 4.155 ;
        RECT  11.550 3.685 12.810 4.155 ;
        RECT  11.205 3.225 11.550 4.155 ;
        RECT  8.350 3.685 11.205 4.155 ;
        RECT  7.990 3.190 8.350 4.155 ;
        RECT  4.735 3.685 7.990 4.155 ;
        RECT  4.395 3.455 4.735 4.155 ;
        RECT  3.675 3.685 4.395 4.155 ;
        RECT  3.335 3.455 3.675 4.155 ;
        RECT  1.250 3.685 3.335 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.580 1.600 13.285 1.940 ;
        RECT  12.350 0.950 12.580 2.760 ;
        RECT  11.615 0.950 12.350 1.180 ;
        RECT  12.060 2.530 12.350 2.760 ;
        RECT  11.875 1.530 12.110 2.300 ;
        RECT  11.270 2.070 11.875 2.300 ;
        RECT  11.385 0.950 11.615 1.830 ;
        RECT  10.690 1.600 11.385 1.830 ;
        RECT  11.040 2.070 11.270 2.995 ;
        RECT  9.775 2.765 11.040 2.995 ;
        RECT  10.235 2.300 10.810 2.530 ;
        RECT  10.235 0.990 10.745 1.220 ;
        RECT  9.120 3.225 10.520 3.455 ;
        RECT  10.005 0.465 10.235 2.530 ;
        RECT  8.570 0.465 10.005 0.695 ;
        RECT  9.545 0.925 9.775 2.995 ;
        RECT  9.040 1.475 9.270 2.500 ;
        RECT  8.890 2.730 9.120 3.455 ;
        RECT  9.030 1.475 9.040 1.705 ;
        RECT  8.930 2.270 9.040 2.500 ;
        RECT  8.800 0.925 9.030 1.705 ;
        RECT  7.645 2.730 8.890 2.960 ;
        RECT  7.885 1.475 8.800 1.705 ;
        RECT  8.340 0.465 8.570 1.245 ;
        RECT  8.215 1.935 8.555 2.470 ;
        RECT  7.495 1.015 8.340 1.245 ;
        RECT  6.920 2.240 8.215 2.470 ;
        RECT  7.545 1.475 7.885 1.890 ;
        RECT  7.415 2.730 7.645 3.250 ;
        RECT  7.265 0.465 7.495 1.245 ;
        RECT  6.285 3.020 7.415 3.250 ;
        RECT  4.875 0.465 7.265 0.695 ;
        RECT  6.870 2.240 6.920 2.650 ;
        RECT  6.640 0.935 6.870 2.650 ;
        RECT  6.055 0.975 6.270 2.630 ;
        RECT  6.040 0.975 6.055 3.210 ;
        RECT  5.860 0.975 6.040 1.210 ;
        RECT  5.825 2.390 6.040 3.210 ;
        RECT  2.675 2.980 5.825 3.210 ;
        RECT  5.555 1.615 5.810 1.955 ;
        RECT  5.325 0.925 5.555 2.750 ;
        RECT  5.220 0.925 5.325 1.265 ;
        RECT  5.210 2.520 5.325 2.750 ;
        RECT  4.940 1.770 5.030 2.110 ;
        RECT  4.710 1.155 4.940 2.740 ;
        RECT  4.645 0.465 4.875 0.925 ;
        RECT  3.765 1.155 4.710 1.385 ;
        RECT  3.835 2.510 4.710 2.740 ;
        RECT  3.230 0.695 4.645 0.925 ;
        RECT  3.000 0.695 3.230 2.270 ;
        RECT  2.445 0.465 2.675 3.210 ;
        RECT  2.060 0.465 2.445 0.695 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFQD0BWP7T

MACRO EDFQD1BWP7T
    CLASS CORE ;
    FOREIGN EDFQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.530 0.470 13.860 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.345 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.100 -0.235 14.000 0.235 ;
        RECT  12.760 -0.235 13.100 0.810 ;
        RECT  11.625 -0.235 12.760 0.235 ;
        RECT  11.395 -0.235 11.625 0.780 ;
        RECT  8.110 -0.235 11.395 0.235 ;
        RECT  7.880 -0.235 8.110 0.785 ;
        RECT  4.415 -0.235 7.880 0.235 ;
        RECT  4.075 -0.235 4.415 0.465 ;
        RECT  3.715 -0.235 4.075 0.235 ;
        RECT  3.375 -0.235 3.715 0.465 ;
        RECT  1.250 -0.235 3.375 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.055 3.685 14.000 4.155 ;
        RECT  12.810 2.240 13.055 4.155 ;
        RECT  11.680 3.685 12.810 4.155 ;
        RECT  11.335 3.225 11.680 4.155 ;
        RECT  8.350 3.685 11.335 4.155 ;
        RECT  7.990 3.190 8.350 4.155 ;
        RECT  4.735 3.685 7.990 4.155 ;
        RECT  4.395 3.455 4.735 4.155 ;
        RECT  3.675 3.685 4.395 4.155 ;
        RECT  3.335 3.455 3.675 4.155 ;
        RECT  1.250 3.685 3.335 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.580 1.600 13.285 1.940 ;
        RECT  12.405 1.020 12.580 2.815 ;
        RECT  12.350 0.550 12.405 2.815 ;
        RECT  12.055 0.550 12.350 1.250 ;
        RECT  12.115 2.565 12.350 3.380 ;
        RECT  11.875 1.530 12.110 2.300 ;
        RECT  11.615 1.020 12.055 1.250 ;
        RECT  11.540 2.070 11.875 2.300 ;
        RECT  11.385 1.020 11.615 1.830 ;
        RECT  11.310 2.070 11.540 2.995 ;
        RECT  10.820 1.600 11.385 1.830 ;
        RECT  9.775 2.765 11.310 2.995 ;
        RECT  10.235 2.300 10.940 2.530 ;
        RECT  10.235 0.990 10.925 1.220 ;
        RECT  9.120 3.225 10.605 3.455 ;
        RECT  10.005 0.465 10.235 2.530 ;
        RECT  8.570 0.465 10.005 0.695 ;
        RECT  9.545 0.925 9.775 2.995 ;
        RECT  9.040 1.475 9.270 2.500 ;
        RECT  8.890 2.730 9.120 3.455 ;
        RECT  9.030 1.475 9.040 1.705 ;
        RECT  8.930 2.270 9.040 2.500 ;
        RECT  8.800 0.925 9.030 1.705 ;
        RECT  7.645 2.730 8.890 2.960 ;
        RECT  7.885 1.475 8.800 1.705 ;
        RECT  8.340 0.465 8.570 1.245 ;
        RECT  8.215 1.935 8.555 2.470 ;
        RECT  7.495 1.015 8.340 1.245 ;
        RECT  6.920 2.240 8.215 2.470 ;
        RECT  7.545 1.475 7.885 1.890 ;
        RECT  7.415 2.730 7.645 3.250 ;
        RECT  7.265 0.465 7.495 1.245 ;
        RECT  6.285 3.020 7.415 3.250 ;
        RECT  4.875 0.465 7.265 0.695 ;
        RECT  6.870 2.240 6.920 2.650 ;
        RECT  6.640 0.935 6.870 2.650 ;
        RECT  6.055 0.975 6.270 2.630 ;
        RECT  6.040 0.975 6.055 3.210 ;
        RECT  5.860 0.975 6.040 1.210 ;
        RECT  5.825 2.390 6.040 3.210 ;
        RECT  2.675 2.980 5.825 3.210 ;
        RECT  5.555 1.615 5.810 1.955 ;
        RECT  5.325 0.925 5.555 2.750 ;
        RECT  5.220 0.925 5.325 1.265 ;
        RECT  5.210 2.520 5.325 2.750 ;
        RECT  4.940 1.770 5.030 2.110 ;
        RECT  4.710 1.155 4.940 2.740 ;
        RECT  4.645 0.465 4.875 0.925 ;
        RECT  3.765 1.155 4.710 1.385 ;
        RECT  3.835 2.510 4.710 2.740 ;
        RECT  3.230 0.695 4.645 0.925 ;
        RECT  3.000 0.695 3.230 2.270 ;
        RECT  2.445 0.465 2.675 3.210 ;
        RECT  2.060 0.465 2.445 0.695 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFQD1BWP7T

MACRO EDFQD2BWP7T
    CLASS CORE ;
    FOREIGN EDFQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.605 1.020 13.860 2.730 ;
        RECT  13.580 0.480 13.605 3.360 ;
        RECT  13.375 0.480 13.580 1.290 ;
        RECT  13.375 2.435 13.580 3.360 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.3915 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 0.980 2.710 ;
        RECT  0.575 2.300 0.700 2.710 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.710 1.585 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.345 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 -0.235 14.560 0.235 ;
        RECT  14.095 -0.235 14.325 1.255 ;
        RECT  12.845 -0.235 14.095 0.235 ;
        RECT  12.615 -0.235 12.845 0.615 ;
        RECT  11.545 -0.235 12.615 0.235 ;
        RECT  11.315 -0.235 11.545 0.535 ;
        RECT  8.110 -0.235 11.315 0.235 ;
        RECT  7.880 -0.235 8.110 0.785 ;
        RECT  4.415 -0.235 7.880 0.235 ;
        RECT  4.075 -0.235 4.415 0.465 ;
        RECT  3.715 -0.235 4.075 0.235 ;
        RECT  3.375 -0.235 3.715 0.465 ;
        RECT  1.250 -0.235 3.375 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 3.685 14.560 4.155 ;
        RECT  14.095 2.255 14.325 4.155 ;
        RECT  12.845 3.685 14.095 4.155 ;
        RECT  12.610 3.250 12.845 4.155 ;
        RECT  11.640 3.685 12.610 4.155 ;
        RECT  11.295 3.250 11.640 4.155 ;
        RECT  8.350 3.685 11.295 4.155 ;
        RECT  7.990 3.190 8.350 4.155 ;
        RECT  4.735 3.685 7.990 4.155 ;
        RECT  4.395 3.455 4.735 4.155 ;
        RECT  3.675 3.685 4.395 4.155 ;
        RECT  3.335 3.455 3.675 4.155 ;
        RECT  1.250 3.685 3.335 4.155 ;
        RECT  0.890 3.190 1.250 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.580 1.600 13.285 1.940 ;
        RECT  12.350 1.020 12.580 2.815 ;
        RECT  11.615 1.020 12.350 1.250 ;
        RECT  12.035 2.585 12.350 2.815 ;
        RECT  11.875 1.600 12.105 2.300 ;
        RECT  11.540 2.070 11.875 2.300 ;
        RECT  11.385 1.020 11.615 1.830 ;
        RECT  11.310 2.070 11.540 2.995 ;
        RECT  10.820 1.600 11.385 1.830 ;
        RECT  9.775 2.765 11.310 2.995 ;
        RECT  10.235 2.300 10.940 2.530 ;
        RECT  10.235 0.990 10.925 1.220 ;
        RECT  9.120 3.225 10.570 3.455 ;
        RECT  10.005 0.465 10.235 2.530 ;
        RECT  8.570 0.465 10.005 0.695 ;
        RECT  9.545 0.925 9.775 2.995 ;
        RECT  9.040 1.475 9.270 2.500 ;
        RECT  8.890 2.730 9.120 3.455 ;
        RECT  9.030 1.475 9.040 1.705 ;
        RECT  8.930 2.270 9.040 2.500 ;
        RECT  8.800 0.925 9.030 1.705 ;
        RECT  7.645 2.730 8.890 2.960 ;
        RECT  7.885 1.475 8.800 1.705 ;
        RECT  8.340 0.465 8.570 1.245 ;
        RECT  8.215 1.935 8.555 2.470 ;
        RECT  7.495 1.015 8.340 1.245 ;
        RECT  6.920 2.240 8.215 2.470 ;
        RECT  7.545 1.475 7.885 1.890 ;
        RECT  7.415 2.730 7.645 3.250 ;
        RECT  7.265 0.465 7.495 1.245 ;
        RECT  6.285 3.020 7.415 3.250 ;
        RECT  4.875 0.465 7.265 0.695 ;
        RECT  6.870 2.240 6.920 2.650 ;
        RECT  6.640 0.935 6.870 2.650 ;
        RECT  6.055 0.975 6.270 2.630 ;
        RECT  6.040 0.975 6.055 3.210 ;
        RECT  5.860 0.975 6.040 1.210 ;
        RECT  5.825 2.390 6.040 3.210 ;
        RECT  2.675 2.980 5.825 3.210 ;
        RECT  5.555 1.615 5.810 1.955 ;
        RECT  5.325 0.925 5.555 2.750 ;
        RECT  5.220 0.925 5.325 1.265 ;
        RECT  5.210 2.520 5.325 2.750 ;
        RECT  4.940 1.770 5.030 2.110 ;
        RECT  4.710 1.155 4.940 2.740 ;
        RECT  4.645 0.465 4.875 0.925 ;
        RECT  3.765 1.155 4.710 1.385 ;
        RECT  3.835 2.510 4.710 2.740 ;
        RECT  3.230 0.695 4.645 0.925 ;
        RECT  3.000 0.695 3.230 2.270 ;
        RECT  2.445 0.465 2.675 3.210 ;
        RECT  2.060 0.465 2.445 0.695 ;
        RECT  2.085 2.815 2.445 3.055 ;
        RECT  1.945 1.205 2.175 2.215 ;
        RECT  0.545 1.205 1.945 1.455 ;
        RECT  0.345 0.635 0.545 1.455 ;
        RECT  0.345 3.065 0.525 3.300 ;
        RECT  0.115 0.635 0.345 3.300 ;
    END
END EDFQD2BWP7T

MACRO FA1D0BWP7T
    CLASS CORE ;
    FOREIGN FA1D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN S
        ANTENNADIFFAREA 0.5962 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.340 1.055 11.620 2.715 ;
        RECT  11.205 1.055 11.340 1.285 ;
        RECT  10.975 2.375 11.340 2.715 ;
        RECT  10.975 0.470 11.205 1.285 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.415 0.470 12.740 2.865 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.3312 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.065 1.210 10.550 1.540 ;
        RECT  9.595 1.210 10.065 1.770 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.4680 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.680 4.340 2.710 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.3708 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.745 0.980 2.150 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.995 -0.235 12.880 0.235 ;
        RECT  11.615 -0.235 11.995 0.675 ;
        RECT  9.800 -0.235 11.615 0.235 ;
        RECT  9.460 -0.235 9.800 0.465 ;
        RECT  4.885 -0.235 9.460 0.235 ;
        RECT  4.655 -0.235 4.885 0.820 ;
        RECT  1.265 -0.235 4.655 0.235 ;
        RECT  0.885 -0.235 1.265 0.785 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.890 3.685 12.880 4.155 ;
        RECT  11.550 3.455 11.890 4.155 ;
        RECT  4.740 3.685 11.550 4.155 ;
        RECT  4.400 3.450 4.740 4.155 ;
        RECT  1.260 3.685 4.400 4.155 ;
        RECT  0.880 3.105 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.935 1.660 12.165 3.225 ;
        RECT  11.205 2.995 11.935 3.225 ;
        RECT  10.975 2.995 11.205 3.455 ;
        RECT  10.745 1.890 11.110 2.120 ;
        RECT  6.925 3.225 10.975 3.455 ;
        RECT  10.515 1.890 10.745 2.995 ;
        RECT  9.040 0.700 10.605 0.930 ;
        RECT  8.275 2.765 10.515 2.995 ;
        RECT  9.040 2.305 10.285 2.535 ;
        RECT  9.040 1.770 9.360 2.000 ;
        RECT  8.810 0.470 9.040 2.535 ;
        RECT  7.745 0.470 8.810 0.700 ;
        RECT  8.275 0.930 8.520 1.160 ;
        RECT  8.045 0.930 8.275 2.995 ;
        RECT  7.555 0.470 7.745 1.845 ;
        RECT  7.515 0.470 7.555 2.615 ;
        RECT  7.325 1.615 7.515 2.615 ;
        RECT  6.925 0.925 7.080 1.155 ;
        RECT  6.695 0.925 6.925 3.455 ;
        RECT  6.605 2.600 6.695 2.940 ;
        RECT  6.075 0.945 6.305 3.220 ;
        RECT  3.780 2.990 6.075 3.220 ;
        RECT  5.565 0.870 5.795 2.540 ;
        RECT  5.375 0.870 5.565 1.305 ;
        RECT  5.160 2.310 5.565 2.540 ;
        RECT  4.845 1.095 5.075 1.945 ;
        RECT  4.425 1.095 4.845 1.325 ;
        RECT  4.195 0.470 4.425 1.325 ;
        RECT  2.505 0.470 4.195 0.700 ;
        RECT  3.780 0.960 3.965 1.300 ;
        RECT  3.550 0.960 3.780 3.220 ;
        RECT  3.225 1.670 3.550 2.010 ;
        RECT  2.975 0.930 3.320 1.160 ;
        RECT  2.975 2.765 3.280 2.995 ;
        RECT  2.735 0.930 2.975 3.455 ;
        RECT  1.720 3.225 2.735 3.455 ;
        RECT  2.275 0.470 2.505 2.910 ;
        RECT  1.490 2.460 1.720 3.455 ;
        RECT  1.440 2.460 1.490 2.690 ;
        RECT  1.210 1.050 1.440 2.690 ;
        RECT  0.465 1.050 1.210 1.280 ;
        RECT  0.465 2.460 1.210 2.690 ;
        RECT  0.235 0.720 0.465 1.280 ;
        RECT  0.235 2.460 0.465 3.385 ;
    END
END FA1D0BWP7T

MACRO FA1D1BWP7T
    CLASS CORE ;
    FOREIGN FA1D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN S
        ANTENNADIFFAREA 0.9720 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.140 1.085 14.420 2.530 ;
        RECT  14.005 1.085 14.140 1.315 ;
        RECT  13.590 2.300 14.140 2.530 ;
        RECT  13.775 0.495 14.005 1.315 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.215 0.495 15.540 2.865 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.6624 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.305 1.210 12.790 1.590 ;
        RECT  11.850 1.210 12.305 1.770 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.4716 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.200 1.680 6.580 2.710 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.465 2.710 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.795 -0.235 15.680 0.235 ;
        RECT  14.415 -0.235 14.795 0.670 ;
        RECT  13.305 -0.235 14.415 0.235 ;
        RECT  13.075 -0.235 13.305 0.850 ;
        RECT  11.880 -0.235 13.075 0.235 ;
        RECT  11.540 -0.235 11.880 0.470 ;
        RECT  7.025 -0.235 11.540 0.235 ;
        RECT  6.795 -0.235 7.025 0.820 ;
        RECT  3.485 -0.235 6.795 0.235 ;
        RECT  3.020 -0.235 3.485 0.465 ;
        RECT  1.980 -0.235 3.020 0.235 ;
        RECT  1.600 -0.235 1.980 1.185 ;
        RECT  0.545 -0.235 1.600 0.235 ;
        RECT  0.165 -0.235 0.545 1.185 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.690 3.685 15.680 4.155 ;
        RECT  14.350 3.220 14.690 4.155 ;
        RECT  6.880 3.685 14.350 4.155 ;
        RECT  6.540 3.450 6.880 4.155 ;
        RECT  3.420 3.685 6.540 4.155 ;
        RECT  3.040 3.250 3.420 4.155 ;
        RECT  1.990 3.685 3.040 4.155 ;
        RECT  1.610 3.250 1.990 4.155 ;
        RECT  0.545 3.685 1.610 4.155 ;
        RECT  0.165 3.070 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.735 1.660 14.965 2.990 ;
        RECT  14.120 2.760 14.735 2.990 ;
        RECT  13.890 2.760 14.120 3.455 ;
        RECT  9.065 3.225 13.890 3.455 ;
        RECT  13.625 1.545 13.855 2.070 ;
        RECT  13.360 1.840 13.625 2.070 ;
        RECT  13.130 1.840 13.360 2.995 ;
        RECT  10.415 2.765 13.130 2.995 ;
        RECT  11.180 0.700 12.685 0.930 ;
        RECT  11.180 2.305 12.525 2.535 ;
        RECT  11.180 1.770 11.500 2.000 ;
        RECT  10.950 0.470 11.180 2.535 ;
        RECT  9.885 0.470 10.950 0.700 ;
        RECT  10.415 0.930 10.660 1.160 ;
        RECT  10.185 0.930 10.415 2.995 ;
        RECT  9.695 0.470 9.885 1.845 ;
        RECT  9.655 0.470 9.695 2.615 ;
        RECT  9.465 1.615 9.655 2.615 ;
        RECT  9.065 0.925 9.220 1.155 ;
        RECT  8.835 0.925 9.065 3.455 ;
        RECT  8.745 2.600 8.835 2.940 ;
        RECT  8.215 0.945 8.445 3.220 ;
        RECT  5.920 2.990 8.215 3.220 ;
        RECT  7.705 0.870 7.935 2.540 ;
        RECT  7.515 0.870 7.705 1.305 ;
        RECT  7.300 2.310 7.705 2.540 ;
        RECT  6.985 1.095 7.215 1.945 ;
        RECT  6.565 1.095 6.985 1.325 ;
        RECT  6.335 0.470 6.565 1.325 ;
        RECT  4.645 0.470 6.335 0.700 ;
        RECT  5.920 0.960 6.105 1.300 ;
        RECT  5.690 0.960 5.920 3.220 ;
        RECT  5.365 1.670 5.690 2.010 ;
        RECT  5.115 0.930 5.460 1.160 ;
        RECT  5.115 2.765 5.420 2.995 ;
        RECT  4.875 0.930 5.115 3.455 ;
        RECT  4.080 3.225 4.875 3.455 ;
        RECT  4.415 0.470 4.645 2.910 ;
        RECT  3.850 2.790 4.080 3.455 ;
        RECT  3.755 1.005 3.985 2.555 ;
        RECT  1.240 2.790 3.850 3.020 ;
        RECT  2.625 1.005 3.755 1.235 ;
        RECT  2.340 2.325 3.755 2.555 ;
        RECT  1.240 1.735 2.915 1.965 ;
        RECT  2.395 0.800 2.625 1.235 ;
        RECT  0.900 0.495 1.240 3.020 ;
    END
END FA1D1BWP7T

MACRO FA1D2BWP7T
    CLASS CORE ;
    FOREIGN FA1D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN S
        ANTENNADIFFAREA 0.9662 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.140 1.085 14.420 2.530 ;
        RECT  13.845 1.085 14.140 1.315 ;
        RECT  13.430 2.300 14.140 2.530 ;
        RECT  13.615 0.945 13.845 1.315 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 0.975 15.540 3.450 ;
        RECT  15.260 0.495 15.285 3.450 ;
        RECT  15.055 0.495 15.260 1.305 ;
        RECT  15.000 3.220 15.260 3.450 ;
        END
    END CO
    PIN CI
        ANTENNAGATEAREA 0.6624 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.690 1.210 13.300 1.590 ;
        RECT  12.410 1.210 12.690 1.825 ;
        END
    END CI
    PIN B
        ANTENNAGATEAREA 0.4716 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.200 1.680 6.580 2.710 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.465 2.710 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.305 ;
        RECT  14.635 -0.235 15.775 0.235 ;
        RECT  14.255 -0.235 14.635 0.670 ;
        RECT  13.155 -0.235 14.255 0.235 ;
        RECT  12.925 -0.235 13.155 0.795 ;
        RECT  11.720 -0.235 12.925 0.235 ;
        RECT  11.430 -0.235 11.720 0.795 ;
        RECT  6.985 -0.235 11.430 0.235 ;
        RECT  6.755 -0.235 6.985 0.820 ;
        RECT  3.485 -0.235 6.755 0.235 ;
        RECT  3.020 -0.235 3.485 0.465 ;
        RECT  1.980 -0.235 3.020 0.235 ;
        RECT  1.600 -0.235 1.980 1.185 ;
        RECT  0.545 -0.235 1.600 0.235 ;
        RECT  0.165 -0.235 0.545 1.185 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.235 16.005 4.155 ;
        RECT  14.530 3.685 15.775 4.155 ;
        RECT  14.190 3.220 14.530 4.155 ;
        RECT  6.880 3.685 14.190 4.155 ;
        RECT  6.540 3.450 6.880 4.155 ;
        RECT  3.420 3.685 6.540 4.155 ;
        RECT  3.040 3.250 3.420 4.155 ;
        RECT  1.990 3.685 3.040 4.155 ;
        RECT  1.610 3.250 1.990 4.155 ;
        RECT  0.545 3.685 1.610 4.155 ;
        RECT  0.165 3.070 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.650 1.660 14.880 2.990 ;
        RECT  13.960 2.760 14.650 2.990 ;
        RECT  13.730 2.760 13.960 3.455 ;
        RECT  13.520 1.725 13.750 2.070 ;
        RECT  9.065 3.225 13.730 3.455 ;
        RECT  13.200 1.840 13.520 2.070 ;
        RECT  12.970 1.840 13.200 2.995 ;
        RECT  10.415 2.765 12.970 2.995 ;
        RECT  12.180 0.700 12.535 0.930 ;
        RECT  11.180 2.305 12.450 2.535 ;
        RECT  11.950 0.700 12.180 1.255 ;
        RECT  11.180 1.025 11.950 1.255 ;
        RECT  11.180 1.770 11.500 2.000 ;
        RECT  10.950 0.470 11.180 2.535 ;
        RECT  9.845 0.470 10.950 0.700 ;
        RECT  10.415 0.930 10.620 1.160 ;
        RECT  10.185 0.930 10.415 2.995 ;
        RECT  9.695 0.470 9.845 1.845 ;
        RECT  9.615 0.470 9.695 2.615 ;
        RECT  9.465 1.615 9.615 2.615 ;
        RECT  9.065 0.925 9.180 1.155 ;
        RECT  8.835 0.925 9.065 3.455 ;
        RECT  8.745 2.600 8.835 2.940 ;
        RECT  8.175 0.945 8.405 3.220 ;
        RECT  5.920 2.990 8.175 3.220 ;
        RECT  7.665 0.870 7.895 2.540 ;
        RECT  7.475 0.870 7.665 1.305 ;
        RECT  7.300 2.310 7.665 2.540 ;
        RECT  6.985 1.095 7.215 1.945 ;
        RECT  6.525 1.095 6.985 1.325 ;
        RECT  6.295 0.470 6.525 1.325 ;
        RECT  4.645 0.470 6.295 0.700 ;
        RECT  5.920 0.960 6.065 1.300 ;
        RECT  5.690 0.960 5.920 3.220 ;
        RECT  5.365 1.670 5.690 2.010 ;
        RECT  5.115 0.930 5.420 1.160 ;
        RECT  5.115 2.765 5.420 2.995 ;
        RECT  4.875 0.930 5.115 3.455 ;
        RECT  4.080 3.225 4.875 3.455 ;
        RECT  4.415 0.470 4.645 2.910 ;
        RECT  3.850 2.790 4.080 3.455 ;
        RECT  3.755 1.005 3.985 2.555 ;
        RECT  1.240 2.790 3.850 3.020 ;
        RECT  2.625 1.005 3.755 1.235 ;
        RECT  2.340 2.325 3.755 2.555 ;
        RECT  1.240 1.735 2.915 1.965 ;
        RECT  2.395 0.800 2.625 1.235 ;
        RECT  0.900 0.495 1.240 3.020 ;
    END
END FA1D2BWP7T

MACRO FILL16BWP7T
    CLASS CORE ;
    FOREIGN FILL16BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 8.960 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 8.960 4.155 ;
        END
    END VDD
END FILL16BWP7T

MACRO FILL1BWP7T
    CLASS CORE ;
    FOREIGN FILL1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 0.560 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 0.560 4.155 ;
        END
    END VDD
END FILL1BWP7T

MACRO FILL2BWP7T
    CLASS CORE ;
    FOREIGN FILL2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 1.120 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 1.120 4.155 ;
        END
    END VDD
END FILL2BWP7T

MACRO FILL32BWP7T
    CLASS CORE ;
    FOREIGN FILL32BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 17.920 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 17.920 4.155 ;
        END
    END VDD
END FILL32BWP7T

MACRO FILL4BWP7T
    CLASS CORE ;
    FOREIGN FILL4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 2.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 2.240 4.155 ;
        END
    END VDD
END FILL4BWP7T

MACRO FILL64BWP7T
    CLASS CORE ;
    FOREIGN FILL64BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 35.840 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 35.840 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 35.840 4.155 ;
        END
    END VDD
END FILL64BWP7T

MACRO FILL8BWP7T
    CLASS CORE ;
    FOREIGN FILL8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 4.480 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 4.480 4.155 ;
        END
    END VDD
END FILL8BWP7T

MACRO GAN2D1BWP7T
    CLASS CORE ;
    FOREIGN GAN2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.180 4.340 2.740 ;
        RECT  2.710 1.180 4.060 1.420 ;
        RECT  2.710 2.500 4.060 2.740 ;
        RECT  2.470 0.640 2.710 1.420 ;
        RECT  2.470 2.500 2.710 3.280 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.715 0.905 2.055 ;
        RECT  0.140 1.715 0.420 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.570 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.930 ;
        RECT  3.550 -0.235 3.940 0.235 ;
        RECT  3.170 -0.235 3.550 0.930 ;
        RECT  0.540 -0.235 3.170 0.235 ;
        RECT  0.160 -0.235 0.540 0.930 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.980 4.320 4.155 ;
        RECT  3.550 3.685 3.940 4.155 ;
        RECT  3.170 2.980 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.990 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.980 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.120 1.715 3.810 2.055 ;
        RECT  1.880 0.690 2.120 2.730 ;
        RECT  1.720 0.690 1.880 0.930 ;
        RECT  1.240 2.490 1.880 2.730 ;
        RECT  0.870 0.465 1.395 0.960 ;
        RECT  1.000 2.490 1.240 3.280 ;
    END
END GAN2D1BWP7T

MACRO GAN2D2BWP7T
    CLASS CORE ;
    FOREIGN GAN2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.180 4.340 2.740 ;
        RECT  3.480 1.180 4.060 1.420 ;
        RECT  3.480 2.500 4.060 2.740 ;
        RECT  3.240 0.640 3.480 1.420 ;
        RECT  3.240 2.500 3.480 3.280 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.715 0.905 2.055 ;
        RECT  0.140 1.715 0.420 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.570 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.930 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.930 ;
        RECT  0.540 -0.235 2.400 0.235 ;
        RECT  0.160 -0.235 0.540 0.930 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.980 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.980 2.780 4.155 ;
        RECT  2.080 3.685 2.400 4.155 ;
        RECT  1.700 2.990 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.980 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.120 1.715 3.810 2.055 ;
        RECT  1.880 0.690 2.120 2.730 ;
        RECT  1.720 0.690 1.880 0.930 ;
        RECT  1.240 2.490 1.880 2.730 ;
        RECT  0.850 0.535 1.360 0.965 ;
        RECT  1.000 2.490 1.240 3.280 ;
    END
END GAN2D2BWP7T

MACRO GAOI21D1BWP7T
    CLASS CORE ;
    FOREIGN GAOI21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 2.3298 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 0.640 4.245 1.390 ;
        RECT  2.705 1.160 4.015 1.390 ;
        RECT  2.660 0.640 2.705 1.390 ;
        RECT  2.380 0.640 2.660 2.680 ;
        RECT  1.775 0.640 2.380 0.980 ;
        RECT  1.235 2.450 2.380 2.680 ;
        RECT  1.005 2.450 1.235 3.280 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.715 3.865 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.715 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 -0.235 4.480 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  0.545 -0.235 3.170 0.235 ;
        RECT  0.165 -0.235 0.545 0.925 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 3.685 4.480 4.155 ;
        RECT  3.175 2.995 3.555 4.155 ;
        RECT  0.000 3.685 3.175 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.870 2.830 4.310 3.365 ;
        RECT  1.715 2.940 2.805 3.225 ;
        RECT  0.870 0.510 1.390 0.960 ;
        RECT  0.170 2.835 0.585 3.390 ;
        LAYER VIA12 ;
        RECT  3.945 2.950 4.205 3.210 ;
        RECT  2.105 2.950 2.365 3.210 ;
        RECT  0.245 2.950 0.505 3.210 ;
        LAYER METAL2 ;
        RECT  0.185 2.940 4.310 3.220 ;
    END
END GAOI21D1BWP7T

MACRO GAOI21D2BWP7T
    CLASS CORE ;
    FOREIGN GAOI21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 3.5996 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.350 0.695 6.580 2.660 ;
        RECT  6.200 0.695 6.350 0.925 ;
        RECT  5.715 2.430 6.350 2.660 ;
        RECT  5.485 2.430 5.715 3.280 ;
        RECT  3.475 2.430 5.485 2.660 ;
        RECT  3.245 2.430 3.475 3.280 ;
        RECT  2.660 2.430 3.245 2.660 ;
        RECT  2.660 0.640 2.760 0.925 ;
        RECT  2.380 0.640 2.660 2.660 ;
        RECT  1.995 0.640 2.380 0.925 ;
        RECT  1.765 0.640 1.995 1.385 ;
        RECT  0.465 1.155 1.765 1.385 ;
        RECT  0.235 0.640 0.465 1.385 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.715 1.625 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.715 5.460 2.150 ;
        RECT  3.810 1.920 5.150 2.150 ;
        RECT  3.500 1.715 3.810 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.210 6.050 2.150 ;
        RECT  3.220 1.210 5.740 1.440 ;
        RECT  2.910 1.210 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.015 -0.235 6.720 0.235 ;
        RECT  4.635 -0.235 5.015 0.925 ;
        RECT  4.320 -0.235 4.635 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  1.310 -0.235 3.940 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 3.685 6.720 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.070 2.890 6.560 3.360 ;
        RECT  5.315 0.525 5.840 0.945 ;
        RECT  4.015 2.940 4.945 3.280 ;
        RECT  3.120 0.485 3.600 0.925 ;
        RECT  2.030 2.940 2.705 3.290 ;
        RECT  1.750 2.405 2.030 3.290 ;
        RECT  0.465 2.405 1.750 2.635 ;
        RECT  0.235 2.405 0.465 3.280 ;
        LAYER VIA12 ;
        RECT  6.240 2.950 6.500 3.210 ;
        RECT  4.335 2.950 4.595 3.210 ;
        RECT  2.105 2.950 2.365 3.210 ;
        LAYER METAL2 ;
        RECT  2.045 2.940 6.560 3.220 ;
    END
END GAOI21D2BWP7T

MACRO GAOI22D1BWP7T
    CLASS CORE ;
    FOREIGN GAOI22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5122 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 2.475 4.245 3.280 ;
        RECT  2.705 2.475 4.015 2.705 ;
        RECT  2.660 0.695 2.760 0.925 ;
        RECT  2.660 2.475 2.705 3.280 ;
        RECT  2.380 0.695 2.660 3.280 ;
        RECT  1.720 0.695 2.380 0.925 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.770 0.980 2.150 ;
        RECT  0.140 1.770 0.420 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.570 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        RECT  3.500 1.770 4.060 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.210 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  0.540 -0.235 3.940 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 3.685 4.480 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.060 2.935 3.665 3.425 ;
        RECT  3.100 0.515 3.620 0.950 ;
        RECT  0.880 0.480 1.355 0.950 ;
        RECT  0.870 2.870 1.355 3.365 ;
        LAYER VIA12 ;
        RECT  3.235 2.950 3.495 3.210 ;
        RECT  0.990 2.945 1.250 3.205 ;
        LAYER METAL2 ;
        RECT  1.310 2.940 3.555 3.220 ;
        RECT  0.930 2.935 1.310 3.220 ;
    END
END GAOI22D1BWP7T

MACRO GBUFFD1BWP7T
    CLASS CORE ;
    FOREIGN GBUFFD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.695 2.100 3.225 ;
        RECT  1.720 0.695 1.820 0.925 ;
        RECT  1.720 2.995 1.820 3.225 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.235 2.240 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 3.685 2.240 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.340 1.155 1.570 2.055 ;
        RECT  0.465 1.155 1.340 1.385 ;
        RECT  0.440 2.995 0.520 3.225 ;
        RECT  0.440 0.640 0.465 1.385 ;
        RECT  0.180 0.640 0.440 3.225 ;
    END
END GBUFFD1BWP7T

MACRO GBUFFD2BWP7T
    CLASS CORE ;
    FOREIGN GBUFFD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.175 4.340 2.710 ;
        RECT  3.475 1.175 4.060 1.405 ;
        RECT  3.475 2.480 4.060 2.710 ;
        RECT  3.245 0.640 3.475 1.405 ;
        RECT  3.245 2.480 3.475 3.280 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.770 1.625 2.000 ;
        RECT  0.140 1.770 0.420 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  2.080 -0.235 2.400 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  2.080 3.685 2.400 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.285 1.715 3.810 2.055 ;
        RECT  2.055 1.170 2.285 2.760 ;
        RECT  1.235 1.170 2.055 1.400 ;
        RECT  1.235 2.530 2.055 2.760 ;
        RECT  1.005 0.640 1.235 1.400 ;
        RECT  1.005 2.530 1.235 3.280 ;
    END
END GBUFFD2BWP7T

MACRO GBUFFD3BWP7T
    CLASS CORE ;
    FOREIGN GBUFFD3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 2.5359 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.725 ;
        RECT  3.475 1.210 4.060 1.445 ;
        RECT  3.475 2.495 4.060 2.725 ;
        RECT  3.245 0.640 3.475 1.445 ;
        RECT  3.245 2.495 3.475 3.280 ;
        RECT  2.005 1.215 3.245 1.445 ;
        RECT  2.005 2.495 3.245 2.725 ;
        RECT  1.775 0.640 2.005 1.445 ;
        RECT  1.775 2.495 2.005 3.280 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.210 0.980 2.165 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.930 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.930 ;
        RECT  1.310 -0.235 2.400 0.235 ;
        RECT  0.930 -0.235 1.310 0.930 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  1.310 3.685 2.400 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.545 1.715 3.810 2.055 ;
        RECT  1.315 1.715 1.545 2.625 ;
        RECT  0.465 2.395 1.315 2.625 ;
        RECT  0.440 0.695 0.520 0.925 ;
        RECT  0.440 2.395 0.465 3.280 ;
        RECT  0.180 0.695 0.440 3.280 ;
    END
END GBUFFD3BWP7T

MACRO GBUFFD8BWP7T
    CLASS CORE ;
    FOREIGN GBUFFD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 5.1192 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  9.690 1.195 10.220 1.475 ;
        RECT  9.690 2.395 10.220 2.675 ;
        RECT  8.790 1.195 9.690 2.675 ;
        RECT  8.280 1.195 8.790 1.475 ;
        RECT  8.280 2.395 8.790 2.675 ;
        END
    END Z
    PIN I
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.715 3.810 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.280 -0.235 13.440 0.235 ;
        RECT  12.900 -0.235 13.280 0.925 ;
        RECT  11.740 -0.235 12.900 0.235 ;
        RECT  11.360 -0.235 11.740 0.925 ;
        RECT  11.040 -0.235 11.360 0.235 ;
        RECT  10.660 -0.235 11.040 0.925 ;
        RECT  9.500 -0.235 10.660 0.235 ;
        RECT  9.120 -0.235 9.500 0.925 ;
        RECT  8.800 -0.235 9.120 0.235 ;
        RECT  8.420 -0.235 8.800 0.925 ;
        RECT  7.260 -0.235 8.420 0.235 ;
        RECT  6.880 -0.235 7.260 0.925 ;
        RECT  6.560 -0.235 6.880 0.235 ;
        RECT  6.180 -0.235 6.560 0.925 ;
        RECT  5.020 -0.235 6.180 0.235 ;
        RECT  4.640 -0.235 5.020 0.925 ;
        RECT  4.320 -0.235 4.640 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  1.310 -0.235 2.400 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.280 3.685 13.440 4.155 ;
        RECT  12.900 2.995 13.280 4.155 ;
        RECT  11.740 3.685 12.900 4.155 ;
        RECT  11.360 2.995 11.740 4.155 ;
        RECT  11.040 3.685 11.360 4.155 ;
        RECT  10.660 2.995 11.040 4.155 ;
        RECT  9.500 3.685 10.660 4.155 ;
        RECT  9.120 2.995 9.500 4.155 ;
        RECT  8.800 3.685 9.120 4.155 ;
        RECT  8.420 2.995 8.800 4.155 ;
        RECT  7.260 3.685 8.420 4.155 ;
        RECT  6.880 2.995 7.260 4.155 ;
        RECT  6.560 3.685 6.880 4.155 ;
        RECT  6.180 2.995 6.560 4.155 ;
        RECT  5.020 3.685 6.180 4.155 ;
        RECT  4.640 2.995 5.020 4.155 ;
        RECT  4.320 3.685 4.640 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  1.310 3.685 2.400 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.915 1.770 12.825 2.000 ;
        RECT  12.205 0.640 12.435 1.510 ;
        RECT  12.205 2.360 12.435 3.280 ;
        RECT  10.195 1.160 12.205 1.510 ;
        RECT  10.195 2.360 12.205 2.710 ;
        RECT  9.965 0.640 10.195 1.510 ;
        RECT  9.965 2.360 10.195 3.280 ;
        RECT  7.955 1.160 9.965 1.510 ;
        RECT  7.955 2.360 9.965 2.710 ;
        RECT  7.725 0.640 7.955 1.510 ;
        RECT  7.725 2.360 7.955 3.280 ;
        RECT  5.715 1.160 7.725 1.510 ;
        RECT  5.715 2.360 7.725 2.710 ;
        RECT  5.485 0.640 5.715 1.510 ;
        RECT  5.485 2.360 5.715 3.280 ;
        RECT  4.685 1.160 4.915 2.760 ;
        RECT  3.475 1.160 4.685 1.390 ;
        RECT  3.475 2.530 4.685 2.760 ;
        RECT  3.245 0.640 3.475 1.390 ;
        RECT  3.245 2.530 3.475 3.280 ;
        RECT  2.005 2.530 3.245 2.760 ;
        RECT  1.775 0.640 2.005 1.390 ;
        RECT  1.775 2.530 2.005 3.280 ;
        RECT  0.465 1.160 1.775 1.390 ;
        RECT  0.465 2.530 1.775 2.760 ;
        RECT  0.440 0.640 0.465 1.390 ;
        RECT  0.440 2.530 0.465 3.280 ;
        RECT  0.210 0.640 0.440 3.280 ;
        LAYER VIA12 ;
        RECT  9.900 1.205 10.160 1.465 ;
        RECT  9.900 2.405 10.160 2.665 ;
        RECT  9.380 1.205 9.640 1.465 ;
        RECT  9.380 2.405 9.640 2.665 ;
        RECT  8.860 1.205 9.120 1.465 ;
        RECT  8.860 2.405 9.120 2.665 ;
        RECT  8.340 1.205 8.600 1.465 ;
        RECT  8.340 2.405 8.600 2.665 ;
    END
END GBUFFD8BWP7T

MACRO GDCAP10BWP7T
    CLASS CORE ;
    FOREIGN GDCAP10BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.470 -0.235 22.400 0.235 ;
        RECT  21.090 -0.235 21.470 0.925 ;
        RECT  20.700 -0.235 21.090 0.235 ;
        RECT  20.320 -0.235 20.700 0.925 ;
        RECT  19.230 -0.235 20.320 0.235 ;
        RECT  18.850 -0.235 19.230 0.925 ;
        RECT  18.460 -0.235 18.850 0.235 ;
        RECT  18.080 -0.235 18.460 0.925 ;
        RECT  16.990 -0.235 18.080 0.235 ;
        RECT  16.610 -0.235 16.990 0.925 ;
        RECT  16.220 -0.235 16.610 0.235 ;
        RECT  15.840 -0.235 16.220 0.925 ;
        RECT  14.750 -0.235 15.840 0.235 ;
        RECT  14.370 -0.235 14.750 0.925 ;
        RECT  13.980 -0.235 14.370 0.235 ;
        RECT  13.600 -0.235 13.980 0.925 ;
        RECT  12.510 -0.235 13.600 0.235 ;
        RECT  12.130 -0.235 12.510 0.925 ;
        RECT  11.740 -0.235 12.130 0.235 ;
        RECT  11.360 -0.235 11.740 0.925 ;
        RECT  10.270 -0.235 11.360 0.235 ;
        RECT  9.890 -0.235 10.270 0.925 ;
        RECT  9.500 -0.235 9.890 0.235 ;
        RECT  9.120 -0.235 9.500 0.925 ;
        RECT  8.030 -0.235 9.120 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  7.260 -0.235 7.650 0.235 ;
        RECT  6.880 -0.235 7.260 0.925 ;
        RECT  5.790 -0.235 6.880 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  5.020 -0.235 5.410 0.235 ;
        RECT  4.640 -0.235 5.020 0.925 ;
        RECT  3.550 -0.235 4.640 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.780 -0.235 3.170 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  1.310 -0.235 2.400 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.540 -0.235 0.930 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.240 3.685 22.400 4.155 ;
        RECT  21.860 2.995 22.240 4.155 ;
        RECT  21.470 3.685 21.860 4.155 ;
        RECT  21.090 2.995 21.470 4.155 ;
        RECT  20.000 3.685 21.090 4.155 ;
        RECT  19.620 2.995 20.000 4.155 ;
        RECT  19.230 3.685 19.620 4.155 ;
        RECT  18.850 2.995 19.230 4.155 ;
        RECT  17.760 3.685 18.850 4.155 ;
        RECT  17.380 2.995 17.760 4.155 ;
        RECT  16.990 3.685 17.380 4.155 ;
        RECT  16.610 2.995 16.990 4.155 ;
        RECT  15.520 3.685 16.610 4.155 ;
        RECT  15.140 2.995 15.520 4.155 ;
        RECT  14.750 3.685 15.140 4.155 ;
        RECT  14.370 2.995 14.750 4.155 ;
        RECT  13.280 3.685 14.370 4.155 ;
        RECT  12.900 2.995 13.280 4.155 ;
        RECT  12.510 3.685 12.900 4.155 ;
        RECT  12.130 2.995 12.510 4.155 ;
        RECT  11.040 3.685 12.130 4.155 ;
        RECT  10.660 2.995 11.040 4.155 ;
        RECT  10.270 3.685 10.660 4.155 ;
        RECT  9.890 2.995 10.270 4.155 ;
        RECT  8.800 3.685 9.890 4.155 ;
        RECT  8.420 2.995 8.800 4.155 ;
        RECT  8.030 3.685 8.420 4.155 ;
        RECT  7.650 2.995 8.030 4.155 ;
        RECT  6.560 3.685 7.650 4.155 ;
        RECT  6.180 2.995 6.560 4.155 ;
        RECT  5.790 3.685 6.180 4.155 ;
        RECT  5.410 2.995 5.790 4.155 ;
        RECT  4.320 3.685 5.410 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  3.550 3.685 3.940 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  1.310 3.685 1.700 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  21.935 0.640 22.165 1.420 ;
        RECT  21.060 1.190 21.935 1.420 ;
        RECT  21.500 1.715 21.730 2.625 ;
        RECT  20.625 2.395 21.500 2.625 ;
        RECT  20.830 1.190 21.060 2.055 ;
        RECT  19.925 1.190 20.830 1.420 ;
        RECT  20.395 2.395 20.625 3.280 ;
        RECT  19.490 2.395 20.395 2.625 ;
        RECT  19.695 0.640 19.925 1.420 ;
        RECT  18.820 1.190 19.695 1.420 ;
        RECT  19.260 1.715 19.490 2.625 ;
        RECT  18.385 2.395 19.260 2.625 ;
        RECT  18.590 1.190 18.820 2.055 ;
        RECT  17.685 1.190 18.590 1.420 ;
        RECT  18.155 2.395 18.385 3.280 ;
        RECT  17.250 2.395 18.155 2.625 ;
        RECT  17.455 0.640 17.685 1.420 ;
        RECT  16.580 1.190 17.455 1.420 ;
        RECT  17.020 1.715 17.250 2.625 ;
        RECT  16.145 2.395 17.020 2.625 ;
        RECT  16.350 1.190 16.580 2.055 ;
        RECT  15.445 1.190 16.350 1.420 ;
        RECT  15.915 2.395 16.145 3.280 ;
        RECT  15.010 2.395 15.915 2.625 ;
        RECT  15.215 0.640 15.445 1.420 ;
        RECT  14.340 1.190 15.215 1.420 ;
        RECT  14.780 1.715 15.010 2.625 ;
        RECT  13.905 2.395 14.780 2.625 ;
        RECT  14.110 1.190 14.340 2.055 ;
        RECT  13.205 1.190 14.110 1.420 ;
        RECT  13.675 2.395 13.905 3.280 ;
        RECT  12.770 2.395 13.675 2.625 ;
        RECT  12.975 0.640 13.205 1.420 ;
        RECT  12.100 1.190 12.975 1.420 ;
        RECT  12.540 1.715 12.770 2.625 ;
        RECT  11.665 2.395 12.540 2.625 ;
        RECT  11.870 1.190 12.100 2.055 ;
        RECT  10.965 1.190 11.870 1.420 ;
        RECT  11.435 2.395 11.665 3.280 ;
        RECT  10.530 2.395 11.435 2.625 ;
        RECT  10.735 0.640 10.965 1.420 ;
        RECT  9.860 1.190 10.735 1.420 ;
        RECT  10.300 1.715 10.530 2.625 ;
        RECT  9.425 2.395 10.300 2.625 ;
        RECT  9.630 1.190 9.860 2.055 ;
        RECT  8.725 1.190 9.630 1.420 ;
        RECT  9.195 2.395 9.425 3.280 ;
        RECT  8.290 2.395 9.195 2.625 ;
        RECT  8.495 0.640 8.725 1.420 ;
        RECT  7.620 1.190 8.495 1.420 ;
        RECT  8.060 1.715 8.290 2.625 ;
        RECT  7.185 2.395 8.060 2.625 ;
        RECT  7.390 1.190 7.620 2.055 ;
        RECT  6.485 1.190 7.390 1.420 ;
        RECT  6.955 2.395 7.185 3.280 ;
        RECT  6.050 2.395 6.955 2.625 ;
        RECT  6.255 0.640 6.485 1.420 ;
        RECT  5.380 1.190 6.255 1.420 ;
        RECT  5.820 1.715 6.050 2.625 ;
        RECT  4.945 2.395 5.820 2.625 ;
        RECT  5.150 1.190 5.380 2.055 ;
        RECT  4.245 1.190 5.150 1.420 ;
        RECT  4.715 2.395 4.945 3.280 ;
        RECT  3.810 2.395 4.715 2.625 ;
        RECT  4.015 0.640 4.245 1.420 ;
        RECT  3.140 1.190 4.015 1.420 ;
        RECT  3.580 1.715 3.810 2.625 ;
        RECT  2.705 2.395 3.580 2.625 ;
        RECT  2.910 1.190 3.140 2.055 ;
        RECT  2.005 1.190 2.910 1.420 ;
        RECT  2.475 2.395 2.705 3.280 ;
        RECT  1.570 2.395 2.475 2.625 ;
        RECT  1.775 0.640 2.005 1.420 ;
        RECT  0.900 1.190 1.775 1.420 ;
        RECT  1.340 1.715 1.570 2.625 ;
        RECT  0.465 2.395 1.340 2.625 ;
        RECT  0.670 1.190 0.900 2.055 ;
        RECT  0.235 2.395 0.465 3.280 ;
    END
END GDCAP10BWP7T

MACRO GDCAP2BWP7T
    CLASS CORE ;
    FOREIGN GDCAP2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 -0.235 4.480 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.780 -0.235 3.170 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  1.310 -0.235 2.400 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.540 -0.235 0.930 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  3.550 3.685 3.940 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  1.310 3.685 1.700 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.015 0.635 4.245 1.465 ;
        RECT  3.140 1.235 4.015 1.465 ;
        RECT  3.580 1.715 3.810 2.600 ;
        RECT  2.705 2.370 3.580 2.600 ;
        RECT  2.910 1.235 3.140 2.055 ;
        RECT  2.005 1.235 2.910 1.465 ;
        RECT  2.475 2.370 2.705 3.280 ;
        RECT  1.570 2.370 2.475 2.600 ;
        RECT  1.775 0.640 2.005 1.465 ;
        RECT  0.900 1.235 1.775 1.465 ;
        RECT  1.340 1.715 1.570 2.600 ;
        RECT  0.465 2.370 1.340 2.600 ;
        RECT  0.670 1.235 0.900 2.055 ;
        RECT  0.235 2.370 0.465 3.280 ;
    END
END GDCAP2BWP7T

MACRO GDCAP3BWP7T
    CLASS CORE ;
    FOREIGN GDCAP3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 -0.235 6.720 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  5.020 -0.235 5.410 0.235 ;
        RECT  4.640 -0.235 5.020 0.925 ;
        RECT  3.550 -0.235 4.640 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.780 -0.235 3.170 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  1.310 -0.235 2.400 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.540 -0.235 0.930 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 3.685 6.720 4.155 ;
        RECT  6.180 2.990 6.560 4.155 ;
        RECT  5.790 3.685 6.180 4.155 ;
        RECT  5.410 2.990 5.790 4.155 ;
        RECT  4.320 3.685 5.410 4.155 ;
        RECT  3.940 2.990 4.320 4.155 ;
        RECT  3.550 3.685 3.940 4.155 ;
        RECT  3.170 2.990 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.990 2.080 4.155 ;
        RECT  1.310 3.685 1.700 4.155 ;
        RECT  0.930 2.990 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.255 0.640 6.485 1.445 ;
        RECT  5.380 1.215 6.255 1.445 ;
        RECT  5.820 1.715 6.050 2.570 ;
        RECT  4.945 2.340 5.820 2.570 ;
        RECT  5.150 1.215 5.380 2.055 ;
        RECT  4.245 1.215 5.150 1.445 ;
        RECT  4.715 2.340 4.945 3.280 ;
        RECT  3.810 2.340 4.715 2.570 ;
        RECT  4.015 0.640 4.245 1.445 ;
        RECT  3.140 1.215 4.015 1.445 ;
        RECT  3.580 1.715 3.810 2.570 ;
        RECT  2.705 2.340 3.580 2.570 ;
        RECT  2.910 1.215 3.140 2.055 ;
        RECT  2.005 1.215 2.910 1.445 ;
        RECT  2.475 2.340 2.705 3.280 ;
        RECT  1.570 2.340 2.475 2.570 ;
        RECT  1.775 0.640 2.005 1.445 ;
        RECT  0.900 1.215 1.775 1.445 ;
        RECT  1.340 1.715 1.570 2.570 ;
        RECT  0.465 2.340 1.340 2.570 ;
        RECT  0.670 1.215 0.900 2.055 ;
        RECT  0.235 2.340 0.465 3.280 ;
    END
END GDCAP3BWP7T

MACRO GDCAP4BWP7T
    CLASS CORE ;
    FOREIGN GDCAP4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 -0.235 8.960 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  7.260 -0.235 7.650 0.235 ;
        RECT  6.880 -0.235 7.260 0.925 ;
        RECT  5.790 -0.235 6.880 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  5.020 -0.235 5.410 0.235 ;
        RECT  4.640 -0.235 5.020 0.925 ;
        RECT  3.550 -0.235 4.640 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.780 -0.235 3.170 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  1.310 -0.235 2.400 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.540 -0.235 0.930 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.800 3.685 8.960 4.155 ;
        RECT  8.420 2.995 8.800 4.155 ;
        RECT  8.030 3.685 8.420 4.155 ;
        RECT  7.650 2.995 8.030 4.155 ;
        RECT  6.560 3.685 7.650 4.155 ;
        RECT  6.180 2.995 6.560 4.155 ;
        RECT  5.790 3.685 6.180 4.155 ;
        RECT  5.410 2.995 5.790 4.155 ;
        RECT  4.320 3.685 5.410 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  3.550 3.685 3.940 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  1.310 3.685 1.700 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.495 0.640 8.725 1.430 ;
        RECT  7.620 1.200 8.495 1.430 ;
        RECT  8.060 1.715 8.290 2.600 ;
        RECT  7.185 2.370 8.060 2.600 ;
        RECT  7.390 1.200 7.620 2.055 ;
        RECT  6.485 1.200 7.390 1.430 ;
        RECT  6.955 2.370 7.185 3.280 ;
        RECT  6.050 2.370 6.955 2.600 ;
        RECT  6.255 0.640 6.485 1.430 ;
        RECT  5.380 1.200 6.255 1.430 ;
        RECT  3.140 1.200 4.015 1.430 ;
        RECT  3.580 1.715 3.810 2.600 ;
        RECT  2.705 2.370 3.580 2.600 ;
        RECT  2.910 1.200 3.140 2.055 ;
        RECT  2.005 1.200 2.910 1.430 ;
        RECT  2.475 2.370 2.705 3.280 ;
        RECT  1.570 2.370 2.475 2.600 ;
        RECT  1.775 0.640 2.005 1.430 ;
        RECT  0.900 1.200 1.775 1.430 ;
        RECT  1.340 1.715 1.570 2.600 ;
        RECT  0.465 2.370 1.340 2.600 ;
        RECT  0.670 1.200 0.900 2.055 ;
        RECT  0.235 2.370 0.465 3.280 ;
        RECT  5.820 1.715 6.050 2.600 ;
        RECT  4.945 2.370 5.820 2.600 ;
        RECT  5.150 1.200 5.380 2.055 ;
        RECT  4.245 1.200 5.150 1.430 ;
        RECT  4.715 2.370 4.945 3.280 ;
        RECT  3.810 2.370 4.715 2.600 ;
        RECT  4.015 0.640 4.245 1.430 ;
    END
END GDCAP4BWP7T

MACRO GDCAPBWP7T
    CLASS CORE ;
    FOREIGN GDCAPBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.235 2.240 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.540 -0.235 0.930 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 3.685 2.240 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  1.310 3.685 1.700 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.775 0.640 2.005 1.425 ;
        RECT  0.900 1.195 1.775 1.425 ;
        RECT  1.340 1.715 1.570 2.745 ;
        RECT  0.465 2.515 1.340 2.745 ;
        RECT  0.670 1.195 0.900 2.055 ;
        RECT  0.235 2.515 0.465 3.280 ;
    END
END GDCAPBWP7T

MACRO GDFCNQD1BWP7T
    CLASS CORE ;
    FOREIGN GDFCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Q
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 0.685 15.540 3.230 ;
        RECT  15.160 0.685 15.260 0.935 ;
        RECT  15.160 2.985 15.260 3.230 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  1.070 1.260 2.150 1.540 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.610 1.820 10.605 2.100 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  12.180 1.260 12.770 1.540 ;
        RECT  11.900 1.260 12.180 2.660 ;
        RECT  5.740 2.380 11.900 2.660 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.750 -0.235 15.680 0.235 ;
        RECT  14.370 -0.235 14.750 0.930 ;
        RECT  11.740 -0.235 14.370 0.235 ;
        RECT  11.360 -0.235 11.740 0.930 ;
        RECT  8.030 -0.235 11.360 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  6.560 -0.235 7.650 0.235 ;
        RECT  6.180 -0.235 6.560 0.930 ;
        RECT  1.310 -0.235 6.180 0.235 ;
        RECT  0.930 -0.235 1.310 0.930 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.750 3.685 15.680 4.155 ;
        RECT  14.370 2.985 14.750 4.155 ;
        RECT  12.490 3.685 14.370 4.155 ;
        RECT  12.150 2.995 12.490 4.155 ;
        RECT  8.010 3.685 12.150 4.155 ;
        RECT  7.670 2.995 8.010 4.155 ;
        RECT  5.790 3.685 7.670 4.155 ;
        RECT  5.410 2.995 5.790 4.155 ;
        RECT  1.310 3.685 5.410 4.155 ;
        RECT  0.930 2.990 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.110 1.715 15.030 2.100 ;
        RECT  13.780 0.685 13.960 0.980 ;
        RECT  13.780 2.890 13.960 3.270 ;
        RECT  13.550 0.685 13.780 3.270 ;
        RECT  13.000 0.685 13.280 3.280 ;
        RECT  12.920 0.685 13.000 0.935 ;
        RECT  12.970 2.450 13.000 3.280 ;
        RECT  11.670 2.450 12.970 2.680 ;
        RECT  12.390 1.260 12.770 2.150 ;
        RECT  12.055 0.530 12.565 1.005 ;
        RECT  11.170 1.715 12.100 2.055 ;
        RECT  11.430 2.450 11.670 3.280 ;
        RECT  10.940 1.210 11.170 2.680 ;
        RECT  10.555 2.910 11.115 3.415 ;
        RECT  10.560 0.510 11.040 0.980 ;
        RECT  10.200 1.210 10.940 1.440 ;
        RECT  10.200 2.450 10.940 2.680 ;
        RECT  10.185 1.705 10.710 2.150 ;
        RECT  9.960 0.640 10.200 1.440 ;
        RECT  9.960 2.450 10.200 3.285 ;
        RECT  8.860 1.770 9.915 2.000 ;
        RECT  9.140 2.870 9.545 3.400 ;
        RECT  9.120 0.640 9.500 1.540 ;
        RECT  8.630 0.685 8.860 3.230 ;
        RECT  8.440 0.685 8.630 0.930 ;
        RECT  8.440 2.990 8.630 3.230 ;
        RECT  7.985 1.665 8.365 2.330 ;
        RECT  7.325 1.210 7.705 2.055 ;
        RECT  7.055 2.915 7.300 3.280 ;
        RECT  7.055 0.685 7.285 0.980 ;
        RECT  6.825 0.685 7.055 3.280 ;
        RECT  6.805 0.685 6.825 1.390 ;
        RECT  5.385 1.160 6.805 1.390 ;
        RECT  6.105 2.890 6.575 3.395 ;
        RECT  5.740 1.630 6.145 2.660 ;
        RECT  5.310 0.475 5.915 0.930 ;
        RECT  5.145 1.160 5.385 2.055 ;
        RECT  4.565 2.870 5.040 3.395 ;
        RECT  3.960 0.685 5.000 0.930 ;
        RECT  4.325 1.175 4.605 2.610 ;
        RECT  3.480 1.175 4.325 1.405 ;
        RECT  3.480 2.380 4.325 2.610 ;
        RECT  3.810 2.890 4.300 3.335 ;
        RECT  3.475 1.675 4.025 2.140 ;
        RECT  3.240 0.640 3.480 1.405 ;
        RECT  3.240 2.380 3.480 3.280 ;
        RECT  2.180 1.770 3.195 2.000 ;
        RECT  1.720 0.685 2.760 0.930 ;
        RECT  2.470 2.295 2.750 3.395 ;
        RECT  1.950 1.770 2.180 2.660 ;
        RECT  1.635 2.940 2.115 3.455 ;
        RECT  0.470 2.420 1.950 2.660 ;
        RECT  1.260 1.210 1.580 2.055 ;
        RECT  0.660 1.340 0.980 2.150 ;
        RECT  0.400 0.690 0.520 0.930 ;
        RECT  0.400 2.420 0.470 3.320 ;
        RECT  0.170 0.690 0.400 3.320 ;
        LAYER VIA12 ;
        RECT  14.440 1.830 14.700 2.090 ;
        RECT  13.640 0.710 13.900 0.970 ;
        RECT  13.590 2.950 13.850 3.210 ;
        RECT  13.010 1.830 13.270 2.090 ;
        RECT  12.450 1.270 12.710 1.530 ;
        RECT  10.755 2.950 11.015 3.210 ;
        RECT  10.720 0.710 10.980 0.970 ;
        RECT  10.285 1.830 10.545 2.090 ;
        RECT  9.225 2.950 9.485 3.210 ;
        RECT  9.180 1.270 9.440 1.530 ;
        RECT  8.045 1.830 8.305 2.090 ;
        RECT  7.385 1.270 7.645 1.530 ;
        RECT  6.970 2.950 7.230 3.210 ;
        RECT  6.900 0.710 7.160 0.970 ;
        RECT  6.220 2.950 6.480 3.210 ;
        RECT  5.815 2.390 6.075 2.650 ;
        RECT  4.675 2.950 4.935 3.210 ;
        RECT  4.335 1.270 4.595 1.530 ;
        RECT  3.980 2.950 4.240 3.210 ;
        RECT  3.570 1.830 3.830 2.090 ;
        RECT  2.480 2.390 2.740 2.650 ;
        RECT  1.790 2.950 2.050 3.210 ;
        RECT  1.290 1.270 1.550 1.530 ;
        RECT  0.670 1.830 0.930 2.090 ;
        LAYER METAL2 ;
        RECT  12.950 1.820 14.760 2.100 ;
        RECT  11.620 0.700 13.960 0.980 ;
        RECT  10.665 2.940 13.910 3.220 ;
        RECT  11.340 0.700 11.620 1.540 ;
        RECT  9.120 1.260 11.340 1.540 ;
        RECT  6.775 0.700 11.060 0.980 ;
        RECT  6.875 2.940 9.560 3.220 ;
        RECT  4.270 1.260 7.705 1.540 ;
        RECT  4.895 2.940 6.540 3.220 ;
        RECT  4.615 2.380 4.895 3.220 ;
        RECT  2.370 2.380 4.615 2.660 ;
        RECT  1.730 2.940 4.335 3.220 ;
    END
END GDFCNQD1BWP7T

MACRO GDFQD1BWP7T
    CLASS CORE ;
    FOREIGN GDFQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Q
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 0.695 13.300 3.225 ;
        RECT  12.920 0.695 13.020 0.925 ;
        RECT  12.920 2.995 13.020 3.225 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.675 1.590 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.510 -0.235 13.440 0.235 ;
        RECT  12.130 -0.235 12.510 0.925 ;
        RECT  10.270 -0.235 12.130 0.235 ;
        RECT  9.890 -0.235 10.270 0.925 ;
        RECT  5.790 -0.235 9.890 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  1.310 -0.235 5.410 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.510 3.685 13.440 4.155 ;
        RECT  12.130 2.995 12.510 4.155 ;
        RECT  10.270 3.685 12.130 4.155 ;
        RECT  9.890 2.995 10.270 4.155 ;
        RECT  5.790 3.685 9.890 4.155 ;
        RECT  5.410 2.995 5.790 4.155 ;
        RECT  1.310 3.685 5.410 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.540 1.175 12.770 2.055 ;
        RECT  11.665 1.175 12.540 1.405 ;
        RECT  11.870 1.715 12.250 2.765 ;
        RECT  11.615 2.995 11.720 3.225 ;
        RECT  11.615 0.640 11.665 1.405 ;
        RECT  11.330 0.640 11.615 3.225 ;
        RECT  10.770 0.695 11.050 3.225 ;
        RECT  10.680 0.695 10.770 0.925 ;
        RECT  10.680 2.995 10.770 3.225 ;
        RECT  10.300 1.715 10.530 2.660 ;
        RECT  9.840 2.380 10.300 2.660 ;
        RECT  9.995 1.210 10.090 1.590 ;
        RECT  9.610 1.210 9.995 2.055 ;
        RECT  8.440 2.995 9.480 3.225 ;
        RECT  9.380 0.640 9.425 0.985 ;
        RECT  9.100 0.640 9.380 1.600 ;
        RECT  8.640 1.210 8.870 2.650 ;
        RECT  8.300 0.590 8.855 0.980 ;
        RECT  7.955 1.210 8.640 1.440 ;
        RECT  7.980 2.420 8.640 2.650 ;
        RECT  7.905 1.670 8.410 2.190 ;
        RECT  7.700 2.420 7.980 3.280 ;
        RECT  7.725 0.640 7.955 1.440 ;
        RECT  7.305 1.770 7.675 2.055 ;
        RECT  6.925 1.770 7.305 2.660 ;
        RECT  6.880 0.615 7.260 1.540 ;
        RECT  6.545 2.995 7.240 3.225 ;
        RECT  6.300 0.695 6.545 3.225 ;
        RECT  6.165 0.695 6.300 0.980 ;
        RECT  6.200 2.420 6.300 3.225 ;
        RECT  5.380 2.420 6.200 2.650 ;
        RECT  5.820 1.190 6.050 2.055 ;
        RECT  4.270 1.190 5.820 1.420 ;
        RECT  5.150 1.715 5.380 2.650 ;
        RECT  4.880 2.940 5.010 3.290 ;
        RECT  3.960 0.695 5.000 0.925 ;
        RECT  4.570 2.305 4.880 3.290 ;
        RECT  3.840 2.895 4.315 3.370 ;
        RECT  4.040 1.190 4.270 2.665 ;
        RECT  3.475 1.190 4.040 1.420 ;
        RECT  3.475 2.435 4.040 2.665 ;
        RECT  3.425 1.650 3.810 2.205 ;
        RECT  3.245 0.640 3.475 1.420 ;
        RECT  3.245 2.435 3.475 3.280 ;
        RECT  2.795 1.770 3.195 2.000 ;
        RECT  2.415 1.160 2.795 2.000 ;
        RECT  2.115 0.695 2.760 0.925 ;
        RECT  2.420 2.310 2.760 3.245 ;
        RECT  1.885 0.695 2.115 3.280 ;
        RECT  1.720 0.695 1.885 0.925 ;
        RECT  1.775 2.890 1.885 3.280 ;
        RECT  0.370 0.695 0.520 0.925 ;
        RECT  0.370 1.160 0.470 1.540 ;
        RECT  0.370 2.925 0.465 3.410 ;
        RECT  0.140 0.695 0.370 3.410 ;
        LAYER VIA12 ;
        RECT  11.930 2.425 12.190 2.685 ;
        RECT  11.345 1.270 11.605 1.530 ;
        RECT  10.780 1.830 11.040 2.090 ;
        RECT  9.950 2.390 10.210 2.650 ;
        RECT  9.770 1.270 10.030 1.530 ;
        RECT  9.110 1.270 9.370 1.530 ;
        RECT  8.475 0.710 8.735 0.970 ;
        RECT  7.995 1.830 8.255 2.090 ;
        RECT  7.710 2.950 7.970 3.210 ;
        RECT  6.985 2.390 7.245 2.650 ;
        RECT  6.940 1.270 7.200 1.530 ;
        RECT  6.225 0.710 6.485 0.970 ;
        RECT  4.590 2.390 4.850 2.650 ;
        RECT  3.975 2.950 4.235 3.210 ;
        RECT  3.435 1.830 3.695 2.090 ;
        RECT  2.475 1.220 2.735 1.480 ;
        RECT  2.475 2.390 2.735 2.650 ;
        RECT  1.845 2.950 2.105 3.210 ;
        RECT  0.200 1.220 0.460 1.480 ;
        RECT  0.150 3.090 0.410 3.350 ;
        LAYER METAL2 ;
        RECT  11.870 2.415 12.250 3.220 ;
        RECT  7.650 2.940 11.870 3.220 ;
        RECT  9.710 1.260 11.665 1.540 ;
        RECT  3.375 1.820 11.100 2.100 ;
        RECT  7.140 2.380 10.280 2.660 ;
        RECT  6.880 1.260 9.430 1.540 ;
        RECT  6.165 0.700 8.795 0.980 ;
        RECT  6.860 2.380 7.140 3.780 ;
        RECT  0.420 3.500 6.860 3.780 ;
        RECT  2.415 2.380 4.910 2.660 ;
        RECT  1.785 2.940 4.295 3.220 ;
        RECT  0.140 1.210 2.795 1.490 ;
        RECT  0.140 3.020 0.420 3.780 ;
    END
END GDFQD1BWP7T

MACRO GFILL10BWP7T
    CLASS CORE ;
    FOREIGN GFILL10BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 22.400 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 22.400 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  21.110 2.995 22.220 3.225 ;
        RECT  21.935 0.640 22.165 1.455 ;
        RECT  21.060 1.225 21.935 1.455 ;
        RECT  21.500 1.715 21.730 2.600 ;
        RECT  20.625 2.370 21.500 2.600 ;
        RECT  20.340 0.695 21.450 0.925 ;
        RECT  20.830 1.225 21.060 2.055 ;
        RECT  19.925 1.225 20.830 1.455 ;
        RECT  20.395 2.370 20.625 3.280 ;
        RECT  19.490 2.370 20.395 2.600 ;
        RECT  18.870 2.995 19.980 3.225 ;
        RECT  19.695 0.640 19.925 1.455 ;
        RECT  18.820 1.225 19.695 1.455 ;
        RECT  19.260 1.715 19.490 2.600 ;
        RECT  18.385 2.370 19.260 2.600 ;
        RECT  18.100 0.695 19.210 0.925 ;
        RECT  18.590 1.225 18.820 2.055 ;
        RECT  17.685 1.225 18.590 1.455 ;
        RECT  18.155 2.370 18.385 3.280 ;
        RECT  17.250 2.370 18.155 2.600 ;
        RECT  16.630 2.995 17.740 3.225 ;
        RECT  17.455 0.640 17.685 1.455 ;
        RECT  16.580 1.225 17.455 1.455 ;
        RECT  17.020 1.715 17.250 2.600 ;
        RECT  16.145 2.370 17.020 2.600 ;
        RECT  15.860 0.695 16.970 0.925 ;
        RECT  16.350 1.225 16.580 2.055 ;
        RECT  15.445 1.225 16.350 1.455 ;
        RECT  15.915 2.370 16.145 3.280 ;
        RECT  15.010 2.370 15.915 2.600 ;
        RECT  14.390 2.995 15.500 3.225 ;
        RECT  15.215 0.640 15.445 1.455 ;
        RECT  14.340 1.225 15.215 1.455 ;
        RECT  14.780 1.715 15.010 2.600 ;
        RECT  13.905 2.370 14.780 2.600 ;
        RECT  13.620 0.695 14.730 0.925 ;
        RECT  14.110 1.225 14.340 2.055 ;
        RECT  13.205 1.225 14.110 1.455 ;
        RECT  13.675 2.370 13.905 3.280 ;
        RECT  12.770 2.370 13.675 2.600 ;
        RECT  12.150 2.995 13.260 3.225 ;
        RECT  12.975 0.640 13.205 1.455 ;
        RECT  12.100 1.225 12.975 1.455 ;
        RECT  12.540 1.715 12.770 2.600 ;
        RECT  11.665 2.370 12.540 2.600 ;
        RECT  11.380 0.695 12.490 0.925 ;
        RECT  11.870 1.225 12.100 2.055 ;
        RECT  10.965 1.225 11.870 1.455 ;
        RECT  11.435 2.370 11.665 3.280 ;
        RECT  10.530 2.370 11.435 2.600 ;
        RECT  9.910 2.995 11.020 3.225 ;
        RECT  10.735 0.640 10.965 1.455 ;
        RECT  9.860 1.225 10.735 1.455 ;
        RECT  10.300 1.715 10.530 2.600 ;
        RECT  9.425 2.370 10.300 2.600 ;
        RECT  9.140 0.695 10.250 0.925 ;
        RECT  9.630 1.225 9.860 2.055 ;
        RECT  8.725 1.225 9.630 1.455 ;
        RECT  9.195 2.370 9.425 3.280 ;
        RECT  8.290 2.370 9.195 2.600 ;
        RECT  7.670 2.995 8.780 3.225 ;
        RECT  8.495 0.640 8.725 1.455 ;
        RECT  7.620 1.225 8.495 1.455 ;
        RECT  8.060 1.715 8.290 2.600 ;
        RECT  7.185 2.370 8.060 2.600 ;
        RECT  6.900 0.695 8.010 0.925 ;
        RECT  7.390 1.225 7.620 2.055 ;
        RECT  6.485 1.225 7.390 1.455 ;
        RECT  6.955 2.370 7.185 3.280 ;
        RECT  6.050 2.370 6.955 2.600 ;
        RECT  5.430 2.995 6.540 3.225 ;
        RECT  6.255 0.640 6.485 1.455 ;
        RECT  5.380 1.225 6.255 1.455 ;
        RECT  5.820 1.715 6.050 2.600 ;
        RECT  4.945 2.370 5.820 2.600 ;
        RECT  4.660 0.695 5.770 0.925 ;
        RECT  5.150 1.225 5.380 2.055 ;
        RECT  4.245 1.225 5.150 1.455 ;
        RECT  4.715 2.370 4.945 3.280 ;
        RECT  3.810 2.370 4.715 2.600 ;
        RECT  3.190 2.995 4.300 3.225 ;
        RECT  4.015 0.640 4.245 1.455 ;
        RECT  3.140 1.225 4.015 1.455 ;
        RECT  3.580 1.715 3.810 2.600 ;
        RECT  2.705 2.370 3.580 2.600 ;
        RECT  2.420 0.695 3.530 0.925 ;
        RECT  2.910 1.225 3.140 2.055 ;
        RECT  2.005 1.225 2.910 1.455 ;
        RECT  2.475 2.370 2.705 3.280 ;
        RECT  1.570 2.370 2.475 2.600 ;
        RECT  0.950 2.995 2.060 3.225 ;
        RECT  1.775 0.640 2.005 1.455 ;
        RECT  0.900 1.225 1.775 1.455 ;
        RECT  1.340 1.715 1.570 2.600 ;
        RECT  0.465 2.370 1.340 2.600 ;
        RECT  0.180 0.695 1.290 0.925 ;
        RECT  0.670 1.225 0.900 2.055 ;
        RECT  0.235 2.370 0.465 3.280 ;
    END
END GFILL10BWP7T

MACRO GFILL2BWP7T
    CLASS CORE ;
    FOREIGN GFILL2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 4.480 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 4.480 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.190 2.995 4.300 3.225 ;
        RECT  4.015 0.640 4.245 1.450 ;
        RECT  3.140 1.220 4.015 1.450 ;
        RECT  3.580 1.715 3.810 2.735 ;
        RECT  2.705 2.505 3.580 2.735 ;
        RECT  2.420 0.695 3.530 0.925 ;
        RECT  2.910 1.220 3.140 2.055 ;
        RECT  2.005 1.220 2.910 1.450 ;
        RECT  2.475 2.505 2.705 3.280 ;
        RECT  1.570 2.505 2.475 2.735 ;
        RECT  0.950 2.995 2.060 3.225 ;
        RECT  1.775 0.640 2.005 1.450 ;
        RECT  0.900 1.220 1.775 1.450 ;
        RECT  1.340 1.715 1.570 2.735 ;
        RECT  0.465 2.505 1.340 2.735 ;
        RECT  0.180 0.695 1.290 0.925 ;
        RECT  0.670 1.220 0.900 2.055 ;
        RECT  0.235 2.505 0.465 3.280 ;
    END
END GFILL2BWP7T

MACRO GFILL3BWP7T
    CLASS CORE ;
    FOREIGN GFILL3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 6.720 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 6.720 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.430 2.995 6.540 3.225 ;
        RECT  6.255 0.640 6.485 1.455 ;
        RECT  5.380 1.225 6.255 1.455 ;
        RECT  5.820 1.715 6.050 2.600 ;
        RECT  4.945 2.370 5.820 2.600 ;
        RECT  4.660 0.695 5.770 0.925 ;
        RECT  5.150 1.225 5.380 2.055 ;
        RECT  4.245 1.225 5.150 1.455 ;
        RECT  4.715 2.370 4.945 3.280 ;
        RECT  3.810 2.370 4.715 2.600 ;
        RECT  3.190 2.995 4.300 3.225 ;
        RECT  4.015 0.640 4.245 1.455 ;
        RECT  3.140 1.225 4.015 1.455 ;
        RECT  3.580 1.715 3.810 2.600 ;
        RECT  2.705 2.370 3.580 2.600 ;
        RECT  2.420 0.695 3.530 0.925 ;
        RECT  2.910 1.225 3.140 2.055 ;
        RECT  2.005 1.225 2.910 1.455 ;
        RECT  2.475 2.370 2.705 3.280 ;
        RECT  1.570 2.370 2.475 2.600 ;
        RECT  0.950 2.995 2.060 3.225 ;
        RECT  1.775 0.640 2.005 1.455 ;
        RECT  0.900 1.225 1.775 1.455 ;
        RECT  1.340 1.715 1.570 2.600 ;
        RECT  0.465 2.370 1.340 2.600 ;
        RECT  0.180 0.695 1.290 0.925 ;
        RECT  0.670 1.225 0.900 2.055 ;
        RECT  0.235 2.370 0.465 3.280 ;
    END
END GFILL3BWP7T

MACRO GFILL4BWP7T
    CLASS CORE ;
    FOREIGN GFILL4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 8.960 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 8.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.670 2.995 8.780 3.225 ;
        RECT  8.495 0.640 8.725 1.455 ;
        RECT  7.620 1.225 8.495 1.455 ;
        RECT  8.060 1.715 8.290 2.600 ;
        RECT  7.185 2.370 8.060 2.600 ;
        RECT  6.900 0.695 8.010 0.925 ;
        RECT  7.390 1.225 7.620 2.055 ;
        RECT  6.485 1.225 7.390 1.455 ;
        RECT  6.955 2.370 7.185 3.280 ;
        RECT  6.050 2.370 6.955 2.600 ;
        RECT  5.430 2.995 6.540 3.225 ;
        RECT  6.255 0.640 6.485 1.455 ;
        RECT  5.380 1.225 6.255 1.455 ;
        RECT  5.820 1.715 6.050 2.600 ;
        RECT  4.945 2.370 5.820 2.600 ;
        RECT  4.660 0.695 5.770 0.925 ;
        RECT  5.150 1.225 5.380 2.055 ;
        RECT  4.245 1.225 5.150 1.455 ;
        RECT  4.715 2.370 4.945 3.280 ;
        RECT  3.810 2.370 4.715 2.600 ;
        RECT  3.190 2.995 4.300 3.225 ;
        RECT  4.015 0.640 4.245 1.455 ;
        RECT  3.140 1.225 4.015 1.455 ;
        RECT  3.580 1.715 3.810 2.600 ;
        RECT  2.705 2.370 3.580 2.600 ;
        RECT  2.420 0.695 3.530 0.925 ;
        RECT  2.910 1.225 3.140 2.055 ;
        RECT  2.005 1.225 2.910 1.455 ;
        RECT  2.475 2.370 2.705 3.280 ;
        RECT  1.570 2.370 2.475 2.600 ;
        RECT  0.950 2.995 2.060 3.225 ;
        RECT  1.775 0.640 2.005 1.455 ;
        RECT  0.900 1.225 1.775 1.455 ;
        RECT  1.340 1.715 1.570 2.600 ;
        RECT  0.465 2.370 1.340 2.600 ;
        RECT  0.180 0.695 1.290 0.925 ;
        RECT  0.670 1.225 0.900 2.055 ;
        RECT  0.235 2.370 0.465 3.280 ;
    END
END GFILL4BWP7T

MACRO GFILLBWP7T
    CLASS CORE ;
    FOREIGN GFILLBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.235 2.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 3.685 2.240 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.950 2.995 2.060 3.225 ;
        RECT  1.775 0.640 2.005 1.465 ;
        RECT  0.900 1.235 1.775 1.465 ;
        RECT  1.340 1.715 1.570 2.680 ;
        RECT  0.465 2.450 1.340 2.680 ;
        RECT  0.180 0.695 1.290 0.925 ;
        RECT  0.670 1.235 0.900 2.055 ;
        RECT  0.235 2.450 0.465 3.280 ;
    END
END GFILLBWP7T

MACRO GINVD1BWP7T
    CLASS CORE ;
    FOREIGN GINVD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 0.695 0.520 0.925 ;
        RECT  0.420 2.995 0.520 3.225 ;
        RECT  0.140 0.695 0.420 3.225 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.715 1.570 2.710 ;
        RECT  0.670 1.715 1.260 2.055 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  1.310 -0.235 1.700 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 3.685 2.240 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  1.310 3.685 1.700 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
END GINVD1BWP7T

MACRO GINVD2BWP7T
    CLASS CORE ;
    FOREIGN GINVD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.155 2.100 2.630 ;
        RECT  1.235 1.155 1.820 1.385 ;
        RECT  1.235 2.400 1.820 2.630 ;
        RECT  1.005 0.640 1.235 1.385 ;
        RECT  1.005 2.400 1.235 3.280 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.715 1.570 2.055 ;
        RECT  0.140 1.715 0.420 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 3.685 2.240 4.155 ;
        RECT  1.705 2.995 2.085 4.155 ;
        RECT  0.540 3.685 1.705 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
END GINVD2BWP7T

MACRO GINVD3BWP7T
    CLASS CORE ;
    FOREIGN GINVD3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5359 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.180 4.340 2.745 ;
        RECT  3.475 1.180 4.060 1.410 ;
        RECT  3.475 2.515 4.060 2.745 ;
        RECT  3.245 0.640 3.475 1.410 ;
        RECT  3.245 2.515 3.475 3.280 ;
        RECT  2.005 1.180 3.245 1.410 ;
        RECT  2.005 2.515 3.245 2.745 ;
        RECT  1.775 0.640 2.005 1.410 ;
        RECT  1.775 2.515 2.005 3.280 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.715 3.810 2.055 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  1.310 -0.235 2.400 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.540 -0.235 0.930 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  1.310 3.685 2.400 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.540 3.685 0.930 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
END GINVD3BWP7T

MACRO GINVD8BWP7T
    CLASS CORE ;
    FOREIGN GINVD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 5.1192 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  4.650 1.260 5.170 1.540 ;
        RECT  4.650 2.380 5.170 2.660 ;
        RECT  3.750 1.260 4.650 2.660 ;
        RECT  3.230 1.260 3.750 1.540 ;
        RECT  3.230 2.380 3.750 2.660 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 3.4128 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.770 8.820 2.710 ;
        RECT  0.615 1.770 8.540 2.000 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.800 -0.235 8.960 0.235 ;
        RECT  8.420 -0.235 8.800 0.925 ;
        RECT  7.260 -0.235 8.420 0.235 ;
        RECT  6.880 -0.235 7.260 0.925 ;
        RECT  6.560 -0.235 6.880 0.235 ;
        RECT  6.180 -0.235 6.560 0.925 ;
        RECT  5.020 -0.235 6.180 0.235 ;
        RECT  4.640 -0.235 5.020 0.925 ;
        RECT  4.320 -0.235 4.640 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  2.080 -0.235 2.400 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.800 3.685 8.960 4.155 ;
        RECT  8.420 2.995 8.800 4.155 ;
        RECT  7.260 3.685 8.420 4.155 ;
        RECT  6.880 2.995 7.260 4.155 ;
        RECT  6.560 3.685 6.880 4.155 ;
        RECT  6.180 2.995 6.560 4.155 ;
        RECT  5.020 3.685 6.180 4.155 ;
        RECT  4.640 2.995 5.020 4.155 ;
        RECT  4.320 3.685 4.640 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  2.080 3.685 2.400 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.725 0.640 7.955 1.540 ;
        RECT  7.725 2.345 7.955 3.280 ;
        RECT  5.715 1.190 7.725 1.540 ;
        RECT  5.715 2.345 7.725 2.695 ;
        RECT  5.485 0.640 5.715 1.540 ;
        RECT  5.485 2.345 5.715 3.280 ;
        RECT  3.475 1.190 5.485 1.540 ;
        RECT  3.475 2.345 5.485 2.695 ;
        RECT  3.245 0.640 3.475 1.540 ;
        RECT  3.245 2.345 3.475 3.280 ;
        RECT  1.235 1.190 3.245 1.540 ;
        RECT  1.235 2.345 3.245 2.695 ;
        RECT  1.005 0.640 1.235 1.540 ;
        RECT  1.005 2.345 1.235 3.280 ;
        LAYER VIA12 ;
        RECT  4.850 2.390 5.110 2.650 ;
        RECT  4.330 1.270 4.590 1.530 ;
        RECT  4.330 2.390 4.590 2.650 ;
        RECT  3.810 1.270 4.070 1.530 ;
        RECT  3.810 2.390 4.070 2.650 ;
        RECT  3.290 1.270 3.550 1.530 ;
        RECT  3.290 2.390 3.550 2.650 ;
        RECT  4.850 1.270 5.110 1.530 ;
    END
END GINVD8BWP7T

MACRO GMUX2D1BWP7T
    CLASS CORE ;
    FOREIGN GMUX2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 0.695 0.520 0.925 ;
        RECT  0.420 2.995 0.520 3.225 ;
        RECT  0.140 0.695 0.420 3.225 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  2.870 1.820 6.075 2.100 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  1.170 1.820 2.150 2.100 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  5.090 2.380 6.070 2.660 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 -0.235 6.720 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  1.310 -0.235 5.410 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 3.685 6.720 4.155 ;
        RECT  5.410 2.995 5.790 4.155 ;
        RECT  1.310 3.685 5.410 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.305 0.640 6.540 3.225 ;
        RECT  6.255 0.640 6.305 1.415 ;
        RECT  6.200 2.995 6.305 3.225 ;
        RECT  3.965 1.185 6.255 1.415 ;
        RECT  5.690 1.660 6.075 2.455 ;
        RECT  5.150 1.715 5.460 2.710 ;
        RECT  4.635 2.940 5.070 3.440 ;
        RECT  3.960 0.695 5.000 0.925 ;
        RECT  3.920 2.365 4.300 3.230 ;
        RECT  3.735 1.185 3.965 2.000 ;
        RECT  3.525 1.770 3.735 2.000 ;
        RECT  3.245 0.640 3.475 1.390 ;
        RECT  3.245 2.375 3.475 3.280 ;
        RECT  2.660 1.660 3.250 2.140 ;
        RECT  2.350 1.160 3.245 1.390 ;
        RECT  2.350 2.375 3.245 2.605 ;
        RECT  2.475 2.885 2.875 3.425 ;
        RECT  1.720 0.695 2.760 0.925 ;
        RECT  2.120 1.160 2.350 2.605 ;
        RECT  1.680 2.940 2.185 3.370 ;
        RECT  0.900 1.160 2.120 1.390 ;
        RECT  1.260 1.715 1.570 2.380 ;
        RECT  0.670 1.160 0.900 2.055 ;
        LAYER VIA12 ;
        RECT  5.755 1.830 6.015 2.090 ;
        RECT  5.175 2.390 5.435 2.650 ;
        RECT  4.715 2.950 4.975 3.210 ;
        RECT  3.980 2.390 4.240 2.650 ;
        RECT  2.930 1.830 3.190 2.090 ;
        RECT  2.555 2.950 2.815 3.210 ;
        RECT  1.860 3.000 2.120 3.260 ;
        RECT  1.285 1.830 1.545 2.090 ;
        LAYER METAL2 ;
        RECT  2.495 2.940 5.035 3.220 ;
        RECT  2.130 2.380 4.300 2.660 ;
        RECT  1.850 2.380 2.130 3.320 ;
    END
END GMUX2D1BWP7T

MACRO GMUX2D2BWP7T
    CLASS CORE ;
    FOREIGN GMUX2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 0.640 1.235 1.460 ;
        RECT  1.005 2.480 1.235 3.280 ;
        RECT  0.420 1.230 1.005 1.460 ;
        RECT  0.420 2.480 1.005 2.710 ;
        RECT  0.140 1.230 0.420 2.710 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  5.040 1.820 8.360 2.100 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.770 3.865 2.100 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  7.320 2.380 8.310 2.660 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 -0.235 8.960 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  3.550 -0.235 7.650 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.080 -0.235 3.170 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 3.685 8.960 4.155 ;
        RECT  7.650 2.995 8.030 4.155 ;
        RECT  3.550 3.685 7.650 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.590 0.640 8.820 3.225 ;
        RECT  8.495 0.640 8.590 1.400 ;
        RECT  8.440 2.995 8.590 3.225 ;
        RECT  6.425 1.170 8.495 1.400 ;
        RECT  7.980 1.645 8.360 2.335 ;
        RECT  7.320 1.715 7.700 2.660 ;
        RECT  6.805 2.890 7.350 3.405 ;
        RECT  6.200 0.695 7.240 0.925 ;
        RECT  6.225 2.330 6.505 3.320 ;
        RECT  6.195 1.170 6.425 2.000 ;
        RECT  5.765 1.770 6.195 2.000 ;
        RECT  5.485 0.640 5.715 1.445 ;
        RECT  5.485 2.405 5.715 3.280 ;
        RECT  4.975 1.675 5.535 2.175 ;
        RECT  4.735 1.215 5.485 1.445 ;
        RECT  4.735 2.405 5.485 2.635 ;
        RECT  4.605 2.890 5.150 3.405 ;
        RECT  3.925 0.695 5.000 0.980 ;
        RECT  4.505 1.215 4.735 2.635 ;
        RECT  1.810 1.215 4.505 1.445 ;
        RECT  3.990 2.330 4.270 3.280 ;
        RECT  2.705 2.485 3.990 2.715 ;
        RECT  2.375 0.465 2.840 0.980 ;
        RECT  2.475 2.485 2.705 3.280 ;
        RECT  1.580 1.215 1.810 2.055 ;
        RECT  0.670 1.715 1.580 2.055 ;
        LAYER VIA12 ;
        RECT  8.040 1.830 8.300 2.090 ;
        RECT  7.380 2.390 7.640 2.650 ;
        RECT  6.900 2.950 7.160 3.210 ;
        RECT  6.235 2.390 6.495 2.650 ;
        RECT  5.100 1.830 5.360 2.090 ;
        RECT  4.695 2.950 4.955 3.210 ;
        RECT  4.000 2.390 4.260 2.650 ;
        RECT  3.985 0.710 4.245 0.970 ;
        RECT  2.460 0.710 2.720 0.970 ;
        LAYER METAL2 ;
        RECT  4.610 2.940 7.225 3.220 ;
        RECT  3.940 2.380 6.555 2.660 ;
        RECT  2.400 0.700 4.305 0.980 ;
    END
END GMUX2D2BWP7T

MACRO GMUX2ND1BWP7T
    CLASS CORE ;
    FOREIGN GMUX2ND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 0.695 0.520 0.925 ;
        RECT  0.420 2.995 0.520 3.225 ;
        RECT  0.140 0.695 0.420 3.225 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  5.065 1.820 8.360 2.100 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.715 3.810 2.150 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  7.240 2.380 8.310 2.660 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 -0.235 8.960 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  3.550 -0.235 7.650 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  1.310 -0.235 3.170 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 3.685 8.960 4.155 ;
        RECT  7.650 2.995 8.030 4.155 ;
        RECT  3.550 3.685 7.650 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  1.310 3.685 3.170 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.590 0.640 8.820 3.225 ;
        RECT  8.495 0.640 8.590 1.395 ;
        RECT  8.440 2.995 8.590 3.225 ;
        RECT  6.180 1.165 8.495 1.395 ;
        RECT  7.980 1.770 8.360 2.595 ;
        RECT  7.320 1.770 7.700 2.660 ;
        RECT  6.845 2.910 7.300 3.380 ;
        RECT  6.200 0.695 7.240 0.925 ;
        RECT  6.175 2.380 6.555 3.225 ;
        RECT  5.950 1.165 6.180 2.000 ;
        RECT  5.765 1.770 5.950 2.000 ;
        RECT  5.485 0.640 5.715 1.410 ;
        RECT  5.485 2.450 5.715 3.280 ;
        RECT  4.945 1.640 5.530 2.220 ;
        RECT  4.670 1.180 5.485 1.410 ;
        RECT  4.670 2.450 5.485 2.680 ;
        RECT  4.660 2.910 5.115 3.380 ;
        RECT  4.190 0.695 5.000 0.925 ;
        RECT  4.440 1.180 4.670 2.680 ;
        RECT  2.565 2.450 4.440 2.680 ;
        RECT  3.845 2.910 4.365 3.455 ;
        RECT  3.960 0.695 4.190 1.400 ;
        RECT  2.705 1.170 3.960 1.400 ;
        RECT  2.330 2.910 2.850 3.450 ;
        RECT  2.475 0.640 2.705 1.400 ;
        RECT  2.335 1.770 2.565 2.680 ;
        RECT  1.285 1.770 2.335 2.000 ;
        RECT  1.775 0.640 2.005 1.435 ;
        RECT  1.775 2.405 2.005 3.280 ;
        RECT  0.900 1.205 1.775 1.435 ;
        RECT  0.900 2.405 1.775 2.635 ;
        RECT  0.670 1.205 0.900 2.635 ;
        LAYER VIA12 ;
        RECT  8.040 1.830 8.300 2.090 ;
        RECT  7.380 2.390 7.640 2.650 ;
        RECT  6.940 2.950 7.200 3.210 ;
        RECT  6.235 2.390 6.495 2.650 ;
        RECT  5.125 1.830 5.385 2.090 ;
        RECT  4.775 2.950 5.035 3.210 ;
        RECT  3.905 2.950 4.165 3.210 ;
        RECT  2.470 2.950 2.730 3.210 ;
        LAYER METAL2 ;
        RECT  4.600 2.940 7.260 3.220 ;
        RECT  4.295 2.380 6.555 2.660 ;
        RECT  3.975 2.380 4.295 3.220 ;
        RECT  2.410 2.940 3.975 3.220 ;
    END
END GMUX2ND1BWP7T

MACRO GMUX2ND2BWP7T
    CLASS CORE ;
    FOREIGN GMUX2ND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 0.640 1.235 1.405 ;
        RECT  1.005 2.535 1.235 3.280 ;
        RECT  0.420 1.175 1.005 1.405 ;
        RECT  0.420 2.535 1.005 2.765 ;
        RECT  0.140 1.175 0.420 2.765 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  5.040 1.820 8.360 2.100 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  3.450 1.820 4.390 2.100 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  7.310 2.380 8.310 2.660 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 -0.235 8.960 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  3.550 -0.235 7.650 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.080 -0.235 3.170 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 3.685 8.960 4.155 ;
        RECT  7.650 2.995 8.030 4.155 ;
        RECT  3.550 3.685 7.650 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.590 0.640 8.820 3.225 ;
        RECT  8.495 0.640 8.590 1.400 ;
        RECT  8.440 2.995 8.590 3.225 ;
        RECT  6.425 1.170 8.495 1.400 ;
        RECT  7.980 1.645 8.360 2.385 ;
        RECT  7.390 1.715 7.700 2.710 ;
        RECT  6.200 0.695 7.240 0.925 ;
        RECT  6.805 2.890 7.240 3.455 ;
        RECT  6.225 2.330 6.505 3.320 ;
        RECT  6.195 1.170 6.425 2.000 ;
        RECT  5.765 1.770 6.195 2.000 ;
        RECT  5.485 0.640 5.715 1.405 ;
        RECT  5.485 2.405 5.715 3.280 ;
        RECT  5.030 1.640 5.535 2.175 ;
        RECT  4.800 1.175 5.485 1.405 ;
        RECT  4.800 2.405 5.485 2.635 ;
        RECT  4.605 2.890 5.105 3.440 ;
        RECT  3.960 0.695 5.000 0.925 ;
        RECT  4.570 1.175 4.800 2.635 ;
        RECT  3.140 1.175 4.570 1.405 ;
        RECT  4.010 2.330 4.340 3.335 ;
        RECT  3.500 1.715 4.055 2.100 ;
        RECT  2.910 1.175 3.140 2.070 ;
        RECT  2.590 0.695 2.760 0.925 ;
        RECT  2.590 2.995 2.760 3.225 ;
        RECT  2.360 0.695 2.590 3.225 ;
        RECT  0.670 1.715 2.360 2.055 ;
        LAYER VIA12 ;
        RECT  8.040 1.830 8.300 2.090 ;
        RECT  7.420 2.390 7.680 2.650 ;
        RECT  6.865 2.950 7.125 3.210 ;
        RECT  6.235 2.390 6.495 2.650 ;
        RECT  5.100 1.830 5.360 2.090 ;
        RECT  4.735 2.950 4.995 3.210 ;
        RECT  4.070 2.390 4.330 2.650 ;
        RECT  3.560 1.830 3.820 2.090 ;
        LAYER METAL2 ;
        RECT  4.675 2.940 7.185 3.220 ;
        RECT  4.010 2.380 6.555 2.660 ;
    END
END GMUX2ND2BWP7T

MACRO GND2D1BWP7T
    CLASS CORE ;
    FOREIGN GND2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2698 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.695 2.100 2.710 ;
        RECT  1.720 0.695 1.820 0.925 ;
        RECT  1.235 2.480 1.820 2.710 ;
        RECT  1.005 2.480 1.235 3.280 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.570 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.770 0.955 2.000 ;
        RECT  0.140 1.770 0.420 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 -0.235 2.240 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 3.685 2.240 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.865 0.480 1.375 0.955 ;
    END
END GND2D1BWP7T

MACRO GND2D2BWP7T
    CLASS CORE ;
    FOREIGN GND2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 3.9644 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  2.030 2.940 4.285 3.220 ;
        LAYER METAL1 ;
        RECT  4.060 0.640 4.340 3.260 ;
        RECT  4.015 0.640 4.060 1.395 ;
        RECT  3.895 2.940 4.060 3.260 ;
        RECT  0.465 1.165 4.015 1.395 ;
        RECT  0.400 2.995 0.520 3.225 ;
        RECT  0.400 0.640 0.465 1.395 ;
        RECT  0.170 0.640 0.400 3.225 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 3.220 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.715 3.810 2.710 ;
        RECT  0.980 2.480 3.500 2.710 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 -0.235 4.480 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  2.080 -0.235 2.400 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.000 -0.235 1.700 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 3.685 4.480 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  1.310 3.685 3.170 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.095 0.485 3.645 0.935 ;
        RECT  1.700 2.940 2.780 3.265 ;
        RECT  0.830 0.485 1.380 0.935 ;
        LAYER VIA12 ;
        RECT  3.955 2.950 4.215 3.210 ;
        RECT  2.095 2.950 2.355 3.210 ;
    END
END GND2D2BWP7T

MACRO GND2D3BWP7T
    CLASS CORE ;
    FOREIGN GND2D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 3.8094 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.140 0.700 2.455 0.980 ;
        LAYER METAL1 ;
        RECT  5.485 2.470 5.715 3.280 ;
        RECT  3.475 2.470 5.485 2.700 ;
        RECT  3.245 2.470 3.475 3.280 ;
        RECT  1.235 2.470 3.245 2.700 ;
        RECT  1.005 2.470 1.235 3.280 ;
        RECT  0.420 2.470 1.005 2.700 ;
        RECT  0.420 0.695 0.520 0.980 ;
        RECT  0.140 0.695 0.420 2.700 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.095 1.715 6.050 2.150 ;
        RECT  3.525 1.715 5.095 2.000 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.630 1.715 3.195 2.000 ;
        RECT  0.670 1.715 1.630 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 -0.235 6.720 0.235 ;
        RECT  6.180 -0.235 6.560 0.925 ;
        RECT  5.020 -0.235 6.180 0.235 ;
        RECT  4.640 -0.235 5.020 0.925 ;
        RECT  4.320 -0.235 4.640 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  0.000 -0.235 3.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 3.685 6.720 4.155 ;
        RECT  6.180 2.995 6.560 4.155 ;
        RECT  5.020 3.685 6.180 4.155 ;
        RECT  4.640 2.995 5.020 4.155 ;
        RECT  4.320 3.685 4.640 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  2.080 3.685 2.400 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.485 0.640 5.715 1.450 ;
        RECT  3.475 1.220 5.485 1.450 ;
        RECT  3.245 0.640 3.475 1.450 ;
        RECT  1.235 1.220 3.245 1.450 ;
        RECT  1.710 0.695 2.760 0.980 ;
        RECT  1.005 0.640 1.235 1.450 ;
        LAYER VIA12 ;
        RECT  2.135 0.710 2.395 0.970 ;
        RECT  0.200 0.710 0.460 0.970 ;
    END
END GND2D3BWP7T

MACRO GND3D1BWP7T
    CLASS CORE ;
    FOREIGN GND3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 2.7220 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 2.445 4.245 3.280 ;
        RECT  2.705 2.445 4.015 2.675 ;
        RECT  2.475 2.445 2.705 3.280 ;
        RECT  1.235 2.445 2.475 2.675 ;
        RECT  1.005 2.445 1.235 3.280 ;
        RECT  0.420 2.445 1.005 2.675 ;
        RECT  0.420 0.695 0.520 0.925 ;
        RECT  0.140 0.695 0.420 2.675 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.665 1.210 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 2.150 ;
        RECT  1.260 1.770 1.820 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.770 3.865 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 -0.235 4.480 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  0.000 -0.235 3.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 3.685 4.480 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.015 0.640 4.245 1.415 ;
        RECT  2.760 1.185 4.015 1.415 ;
        RECT  2.530 0.695 2.760 1.415 ;
        RECT  1.720 0.695 2.530 0.925 ;
        RECT  0.805 0.500 1.420 0.950 ;
    END
END GND3D1BWP7T

MACRO GND3D2BWP7T
    CLASS CORE ;
    FOREIGN GND3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 3.2794 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL2 ;
        RECT  0.930 2.940 5.790 3.220 ;
        LAYER METAL1 ;
        RECT  0.980 2.505 1.260 3.280 ;
        RECT  0.420 2.505 0.980 2.735 ;
        RECT  0.420 0.695 0.520 0.925 ;
        RECT  0.140 0.695 0.420 2.735 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.770 3.865 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.225 1.770 5.460 2.150 ;
        RECT  4.995 1.770 5.225 2.610 ;
        RECT  1.750 2.380 4.995 2.610 ;
        RECT  1.520 1.770 1.750 2.610 ;
        RECT  1.260 1.770 1.520 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.210 6.050 2.150 ;
        RECT  0.980 1.210 5.740 1.440 ;
        RECT  0.670 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 -0.235 6.720 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  0.000 -0.235 3.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 3.685 6.720 4.155 ;
        RECT  6.180 2.995 6.560 4.155 ;
        RECT  5.020 3.685 6.180 4.155 ;
        RECT  4.640 2.995 5.020 4.155 ;
        RECT  4.320 3.685 4.640 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  2.080 3.685 2.400 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.345 0.695 6.575 2.765 ;
        RECT  6.200 0.695 6.345 0.925 ;
        RECT  5.740 2.535 6.345 2.765 ;
        RECT  5.310 0.475 5.870 0.965 ;
        RECT  5.460 2.535 5.740 3.280 ;
        RECT  3.960 0.695 5.000 0.925 ;
        RECT  3.135 2.845 3.585 3.440 ;
        RECT  1.720 0.695 2.760 0.925 ;
        RECT  0.820 0.530 1.440 0.975 ;
        LAYER VIA12 ;
        RECT  5.470 2.950 5.730 3.210 ;
        RECT  3.230 2.950 3.490 3.210 ;
        RECT  0.990 2.950 1.250 3.210 ;
    END
END GND3D2BWP7T

MACRO GNR2D1BWP7T
    CLASS CORE ;
    FOREIGN GNR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2661 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.180 2.100 3.225 ;
        RECT  1.235 1.180 1.820 1.410 ;
        RECT  1.720 2.995 1.820 3.225 ;
        RECT  1.005 0.640 1.235 1.410 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.715 1.570 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.770 0.955 2.000 ;
        RECT  0.140 1.770 0.420 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 3.685 2.240 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.830 2.945 1.410 3.440 ;
    END
END GNR2D1BWP7T

MACRO GNR2D2BWP7T
    CLASS CORE ;
    FOREIGN GNR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5322 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.160 4.340 3.225 ;
        RECT  3.475 1.160 4.060 1.390 ;
        RECT  3.960 2.995 4.060 3.225 ;
        RECT  3.245 0.640 3.475 1.390 ;
        RECT  1.235 1.160 3.245 1.390 ;
        RECT  1.005 0.640 1.235 1.390 ;
        RECT  0.375 1.160 1.005 1.390 ;
        RECT  0.375 2.995 0.520 3.225 ;
        RECT  0.145 1.160 0.375 3.225 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.715 3.810 2.660 ;
        RECT  0.980 2.430 3.500 2.660 ;
        RECT  0.670 1.715 0.980 2.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  2.080 -0.235 2.400 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 3.685 4.480 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  2.080 3.685 2.400 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.000 3.685 1.700 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.070 2.935 3.635 3.440 ;
        RECT  0.830 2.935 1.395 3.440 ;
    END
END GNR2D2BWP7T

MACRO GNR3D1BWP7T
    CLASS CORE ;
    FOREIGN GNR3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8061 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.245 0.640 3.475 1.400 ;
        RECT  1.235 1.170 3.245 1.400 ;
        RECT  1.005 0.640 1.235 1.400 ;
        RECT  0.420 1.170 1.005 1.400 ;
        RECT  0.420 2.995 0.520 3.225 ;
        RECT  0.140 1.170 0.420 3.225 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.770 4.340 2.710 ;
        RECT  2.855 1.770 4.060 2.000 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.715 1.570 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  2.080 -0.235 2.400 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.780 3.685 3.940 4.155 ;
        RECT  2.400 2.995 2.780 4.155 ;
        RECT  0.000 3.685 2.400 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.245 2.525 3.475 3.280 ;
        RECT  2.095 2.525 3.245 2.755 ;
        RECT  1.865 2.525 2.095 3.225 ;
        RECT  1.720 2.995 1.865 3.225 ;
        RECT  0.835 2.965 1.390 3.430 ;
    END
END GNR3D1BWP7T

MACRO GNR3D2BWP7T
    CLASS CORE ;
    FOREIGN GNR3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0722 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.485 0.640 5.715 1.395 ;
        RECT  3.475 1.165 5.485 1.395 ;
        RECT  3.245 0.640 3.475 1.395 ;
        RECT  2.100 1.165 3.245 1.395 ;
        RECT  1.820 1.165 2.100 3.280 ;
        RECT  1.235 1.165 1.820 1.395 ;
        RECT  1.775 2.480 1.820 3.280 ;
        RECT  0.465 2.480 1.775 2.710 ;
        RECT  1.005 0.640 1.235 1.395 ;
        RECT  0.235 2.480 0.465 3.280 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.770 6.580 2.710 ;
        RECT  5.095 1.770 6.300 2.000 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.770 3.940 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.570 1.715 1.570 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 -0.235 6.720 0.235 ;
        RECT  6.180 -0.235 6.560 0.925 ;
        RECT  5.020 -0.235 6.180 0.235 ;
        RECT  4.640 -0.235 5.020 0.925 ;
        RECT  4.320 -0.235 4.640 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  2.780 -0.235 3.940 0.235 ;
        RECT  2.400 -0.235 2.780 0.925 ;
        RECT  2.080 -0.235 2.400 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 3.685 6.720 4.155 ;
        RECT  6.180 2.995 6.560 4.155 ;
        RECT  5.020 3.685 6.180 4.155 ;
        RECT  4.640 2.995 5.020 4.155 ;
        RECT  0.000 3.685 4.640 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.485 2.435 5.715 3.280 ;
        RECT  3.475 2.435 5.485 2.665 ;
        RECT  3.875 2.940 4.375 3.425 ;
        RECT  3.245 2.435 3.475 3.280 ;
        RECT  2.345 2.940 2.825 3.425 ;
        RECT  0.875 2.940 1.355 3.425 ;
        LAYER VIA12 ;
        RECT  3.980 2.950 4.240 3.210 ;
        RECT  2.460 2.950 2.720 3.210 ;
        RECT  0.990 2.950 1.250 3.210 ;
        LAYER METAL2 ;
        RECT  0.895 2.940 4.390 3.220 ;
    END
END GNR3D2BWP7T

MACRO GOAI21D1BWP7T
    CLASS CORE ;
    FOREIGN GOAI21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 3.2383 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 2.400 4.245 3.280 ;
        RECT  2.765 2.400 4.015 2.630 ;
        RECT  2.660 2.400 2.765 3.225 ;
        RECT  2.380 1.210 2.660 3.225 ;
        RECT  2.005 1.210 2.380 1.440 ;
        RECT  1.720 2.995 2.380 3.225 ;
        RECT  1.775 0.640 2.005 1.440 ;
        RECT  0.465 1.210 1.775 1.440 ;
        RECT  0.235 0.640 0.465 1.440 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.715 3.930 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.715 1.570 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 -0.235 4.480 0.235 ;
        RECT  3.145 -0.235 3.555 0.925 ;
        RECT  0.000 -0.235 3.145 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 3.685 4.480 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  0.545 3.685 3.170 4.155 ;
        RECT  0.165 2.995 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.840 0.520 4.300 1.015 ;
        RECT  2.300 0.520 2.830 0.980 ;
        RECT  0.865 2.960 1.415 3.445 ;
        RECT  0.860 0.520 1.390 0.980 ;
        LAYER VIA12 ;
        RECT  3.950 0.710 4.210 0.970 ;
        RECT  2.430 0.710 2.690 0.970 ;
        RECT  0.990 0.710 1.250 0.970 ;
        LAYER METAL2 ;
        RECT  0.925 0.700 4.305 0.980 ;
    END
END GOAI21D1BWP7T

MACRO GOAI21D2BWP7T
    CLASS CORE ;
    FOREIGN GOAI21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 4.3120 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.280 0.695 6.540 3.280 ;
        RECT  6.200 0.695 6.280 0.925 ;
        RECT  5.000 1.210 6.280 1.440 ;
        RECT  6.255 2.440 6.280 3.280 ;
        RECT  4.660 0.695 5.000 1.440 ;
        RECT  4.300 1.210 4.660 1.440 ;
        RECT  3.955 0.695 4.300 1.440 ;
        RECT  2.760 1.210 3.955 1.440 ;
        RECT  2.660 0.695 2.760 1.440 ;
        RECT  2.660 2.380 2.710 3.280 ;
        RECT  2.475 0.695 2.660 3.280 ;
        RECT  2.380 0.695 2.475 2.670 ;
        RECT  1.235 2.380 2.380 2.670 ;
        RECT  1.005 2.380 1.235 3.280 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.770 1.625 2.000 ;
        RECT  0.140 1.770 0.420 2.710 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 5.460 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.920 1.670 6.050 2.150 ;
        RECT  5.690 1.670 5.920 2.660 ;
        RECT  3.220 2.380 5.690 2.660 ;
        RECT  2.975 1.670 3.220 2.660 ;
        RECT  2.910 1.670 2.975 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 -0.235 6.720 0.235 ;
        RECT  1.705 -0.235 2.085 0.925 ;
        RECT  0.540 -0.235 1.705 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 3.685 6.720 4.155 ;
        RECT  4.640 2.995 5.020 4.155 ;
        RECT  4.320 3.685 4.640 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  2.080 3.685 3.940 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.320 2.945 5.890 3.425 ;
        RECT  5.355 0.535 5.825 0.980 ;
        RECT  3.080 2.945 3.650 3.425 ;
        RECT  3.110 0.535 3.580 0.980 ;
        RECT  0.850 0.570 1.395 0.980 ;
        LAYER VIA12 ;
        RECT  5.470 0.710 5.730 0.970 ;
        RECT  3.205 0.710 3.465 0.970 ;
        RECT  0.985 0.710 1.245 0.970 ;
        LAYER METAL2 ;
        RECT  0.910 0.700 5.790 0.980 ;
    END
END GOAI21D2BWP7T

MACRO GOR2D1BWP7T
    CLASS CORE ;
    FOREIGN GOR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.165 4.340 2.670 ;
        RECT  2.705 1.165 4.060 1.395 ;
        RECT  2.705 2.440 4.060 2.670 ;
        RECT  2.475 0.640 2.705 1.395 ;
        RECT  2.475 2.440 2.705 3.280 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.715 1.570 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.925 ;
        RECT  3.550 -0.235 3.940 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.080 -0.235 3.170 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.995 4.320 4.155 ;
        RECT  3.550 3.685 3.940 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  0.540 3.685 3.170 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.100 1.715 3.810 2.055 ;
        RECT  1.870 1.225 2.100 3.225 ;
        RECT  1.235 1.225 1.870 1.455 ;
        RECT  1.720 2.995 1.870 3.225 ;
        RECT  0.840 2.965 1.445 3.400 ;
        RECT  1.005 0.640 1.235 1.455 ;
    END
END GOR2D1BWP7T

MACRO GOR2D2BWP7T
    CLASS CORE ;
    FOREIGN GOR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 2.5122 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.640 4.340 3.280 ;
        RECT  4.015 0.640 4.060 1.395 ;
        RECT  4.015 2.440 4.060 3.280 ;
        RECT  2.705 1.165 4.015 1.395 ;
        RECT  2.705 2.440 4.015 2.670 ;
        RECT  2.475 0.640 2.705 1.395 ;
        RECT  2.475 2.440 2.705 3.280 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.715 0.980 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.715 1.570 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 -0.235 4.480 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.080 -0.235 3.170 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 3.685 4.480 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  0.540 3.685 3.170 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.100 1.715 3.810 2.055 ;
        RECT  1.870 1.225 2.100 3.225 ;
        RECT  1.235 1.225 1.870 1.455 ;
        RECT  1.720 2.995 1.870 3.225 ;
        RECT  0.865 2.950 1.395 3.425 ;
        RECT  1.005 0.640 1.235 1.455 ;
    END
END GOR2D2BWP7T

MACRO GSDFCNQD1BWP7T
    CLASS CORE ;
    FOREIGN GSDFCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN SI
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.770 0.955 2.000 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  1.260 1.260 3.195 1.540 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.740 0.685 20.020 3.230 ;
        RECT  19.640 0.685 19.740 0.935 ;
        RECT  19.640 2.985 19.740 3.230 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.210 5.460 2.235 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  5.790 1.820 15.085 2.100 ;
        LAYER METAL1 ;
        RECT  5.740 1.210 6.120 2.150 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  16.940 0.140 17.220 1.600 ;
        RECT  10.500 0.140 16.940 0.420 ;
        RECT  10.500 1.260 10.625 1.540 ;
        RECT  10.220 0.140 10.500 1.540 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.230 -0.235 20.160 0.235 ;
        RECT  18.850 -0.235 19.230 0.930 ;
        RECT  16.220 -0.235 18.850 0.235 ;
        RECT  15.840 -0.235 16.220 0.930 ;
        RECT  12.510 -0.235 15.840 0.235 ;
        RECT  12.130 -0.235 12.510 0.925 ;
        RECT  11.040 -0.235 12.130 0.235 ;
        RECT  10.660 -0.235 11.040 0.930 ;
        RECT  5.790 -0.235 10.660 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  1.295 -0.235 5.410 0.235 ;
        RECT  0.915 -0.235 1.295 0.945 ;
        RECT  0.000 -0.235 0.915 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.230 3.685 20.160 4.155 ;
        RECT  18.850 2.985 19.230 4.155 ;
        RECT  16.970 3.685 18.850 4.155 ;
        RECT  16.630 2.995 16.970 4.155 ;
        RECT  12.490 3.685 16.630 4.155 ;
        RECT  12.150 2.995 12.490 4.155 ;
        RECT  10.270 3.685 12.150 4.155 ;
        RECT  9.890 2.980 10.270 4.155 ;
        RECT  5.790 3.685 9.890 4.155 ;
        RECT  5.410 2.990 5.790 4.155 ;
        RECT  1.295 3.685 5.410 4.155 ;
        RECT  0.950 2.990 1.295 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.590 1.715 19.510 2.100 ;
        RECT  18.260 0.685 18.440 0.980 ;
        RECT  18.260 2.890 18.440 3.280 ;
        RECT  18.030 0.685 18.260 3.280 ;
        RECT  17.480 0.685 17.760 3.280 ;
        RECT  17.400 0.685 17.480 0.935 ;
        RECT  17.450 2.450 17.480 3.280 ;
        RECT  16.150 2.450 17.450 2.680 ;
        RECT  16.905 1.185 17.250 2.150 ;
        RECT  16.505 0.465 17.085 0.930 ;
        RECT  15.650 1.715 16.580 2.055 ;
        RECT  15.910 2.450 16.150 3.280 ;
        RECT  15.420 1.210 15.650 2.680 ;
        RECT  15.110 0.465 15.550 0.980 ;
        RECT  15.130 2.920 15.545 3.435 ;
        RECT  14.680 1.210 15.420 1.440 ;
        RECT  14.680 2.450 15.420 2.680 ;
        RECT  14.665 1.705 15.190 2.150 ;
        RECT  14.440 0.640 14.680 1.440 ;
        RECT  14.440 2.450 14.680 3.285 ;
        RECT  13.340 1.770 14.395 2.000 ;
        RECT  13.930 1.260 14.035 1.540 ;
        RECT  13.615 2.870 14.000 3.435 ;
        RECT  13.655 0.640 13.930 1.540 ;
        RECT  13.110 0.685 13.340 3.230 ;
        RECT  12.920 0.685 13.110 0.930 ;
        RECT  12.920 2.990 13.110 3.230 ;
        RECT  12.465 1.665 12.845 2.330 ;
        RECT  11.805 1.745 12.185 2.660 ;
        RECT  11.535 2.940 11.790 3.280 ;
        RECT  11.535 0.685 11.720 0.980 ;
        RECT  11.305 0.685 11.535 3.280 ;
        RECT  11.285 0.685 11.305 2.630 ;
        RECT  9.865 2.400 11.285 2.630 ;
        RECT  10.640 2.870 11.025 3.435 ;
        RECT  10.220 1.210 10.625 2.055 ;
        RECT  9.835 0.510 10.350 0.980 ;
        RECT  9.625 1.715 9.865 2.630 ;
        RECT  9.150 2.870 9.535 3.435 ;
        RECT  8.440 0.685 9.480 0.930 ;
        RECT  8.805 1.175 9.035 2.660 ;
        RECT  8.325 2.890 8.840 3.415 ;
        RECT  7.960 1.175 8.805 1.405 ;
        RECT  7.960 2.380 8.805 2.660 ;
        RECT  7.955 1.675 8.505 2.140 ;
        RECT  7.720 0.640 7.960 1.405 ;
        RECT  7.720 2.380 7.960 3.280 ;
        RECT  6.720 1.765 7.675 2.005 ;
        RECT  6.950 0.465 7.335 1.030 ;
        RECT  6.950 2.870 7.335 3.435 ;
        RECT  6.490 0.695 6.720 3.225 ;
        RECT  6.200 0.695 6.490 0.925 ;
        RECT  6.200 2.995 6.490 3.225 ;
        RECT  4.830 0.690 5.000 0.930 ;
        RECT  4.830 2.995 5.000 3.230 ;
        RECT  4.550 0.690 4.830 3.230 ;
        RECT  3.960 0.690 4.550 0.930 ;
        RECT  4.040 1.685 4.320 3.280 ;
        RECT  4.010 2.935 4.040 3.280 ;
        RECT  3.580 1.710 3.810 2.460 ;
        RECT  2.995 2.940 3.700 3.280 ;
        RECT  2.220 2.230 3.580 2.460 ;
        RECT  3.160 0.465 3.545 1.030 ;
        RECT  2.780 1.260 3.195 2.000 ;
        RECT  2.450 0.500 2.875 1.030 ;
        RECT  2.450 2.690 2.740 3.405 ;
        RECT  1.990 0.695 2.220 3.225 ;
        RECT  1.720 0.695 1.990 0.925 ;
        RECT  1.720 2.995 1.990 3.225 ;
        RECT  1.260 1.260 1.640 2.175 ;
        RECT  0.120 0.465 0.585 0.980 ;
        RECT  0.185 2.645 0.465 3.435 ;
        LAYER VIA12 ;
        RECT  18.920 1.830 19.180 2.090 ;
        RECT  18.120 2.950 18.380 3.210 ;
        RECT  17.490 1.830 17.750 2.090 ;
        RECT  16.950 1.270 17.210 1.530 ;
        RECT  15.205 0.710 15.465 0.970 ;
        RECT  15.195 2.950 15.455 3.210 ;
        RECT  14.765 1.830 15.025 2.090 ;
        RECT  13.715 1.270 13.975 1.530 ;
        RECT  13.645 2.950 13.905 3.210 ;
        RECT  12.525 1.830 12.785 2.090 ;
        RECT  11.865 2.390 12.125 2.650 ;
        RECT  11.435 2.950 11.695 3.210 ;
        RECT  11.355 0.710 11.615 0.970 ;
        RECT  10.700 2.950 10.960 3.210 ;
        RECT  10.295 1.270 10.555 1.530 ;
        RECT  9.245 2.950 9.505 3.210 ;
        RECT  8.710 2.390 8.970 2.650 ;
        RECT  8.480 2.950 8.740 3.210 ;
        RECT  8.050 1.830 8.310 2.090 ;
        RECT  7.015 2.950 7.275 3.210 ;
        RECT  6.960 0.660 7.220 0.920 ;
        RECT  5.850 1.830 6.110 2.090 ;
        RECT  4.560 2.390 4.820 2.650 ;
        RECT  4.050 1.830 4.310 2.090 ;
        RECT  3.230 2.950 3.490 3.210 ;
        RECT  3.225 0.660 3.485 0.920 ;
        RECT  2.840 1.270 3.100 1.530 ;
        RECT  2.465 2.950 2.725 3.210 ;
        RECT  2.460 0.660 2.720 0.920 ;
        RECT  1.320 1.270 1.580 1.530 ;
        RECT  0.235 0.660 0.495 0.920 ;
        RECT  0.195 2.950 0.455 3.210 ;
        LAYER METAL2 ;
        RECT  17.430 1.820 19.240 2.100 ;
        RECT  16.045 2.940 18.440 3.220 ;
        RECT  15.765 1.260 16.045 3.220 ;
        RECT  13.625 1.260 15.765 1.540 ;
        RECT  15.100 2.940 15.765 3.220 ;
        RECT  11.270 0.700 15.560 0.980 ;
        RECT  11.325 2.940 13.965 3.220 ;
        RECT  8.640 2.380 12.215 2.660 ;
        RECT  9.465 2.940 11.030 3.220 ;
        RECT  9.185 2.940 9.465 3.780 ;
        RECT  7.505 3.500 9.185 3.780 ;
        RECT  8.085 2.940 8.825 3.220 ;
        RECT  7.805 2.380 8.085 3.220 ;
        RECT  6.020 2.380 7.805 2.660 ;
        RECT  7.225 2.940 7.505 3.780 ;
        RECT  3.165 0.650 7.285 0.930 ;
        RECT  6.925 2.940 7.225 3.220 ;
        RECT  5.740 2.380 6.020 3.220 ;
        RECT  3.170 2.940 5.740 3.220 ;
        RECT  2.735 2.380 4.880 2.660 ;
        RECT  1.770 1.820 4.375 2.100 ;
        RECT  0.175 0.650 2.780 0.930 ;
        RECT  2.450 2.380 2.735 3.285 ;
        RECT  1.490 1.820 1.770 2.710 ;
        RECT  0.465 2.430 1.490 2.710 ;
        RECT  0.185 2.430 0.465 3.270 ;
    END
END GSDFCNQD1BWP7T

MACRO GTIEHBWP7T
    CLASS CORE ;
    FOREIGN GTIEHBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 0.7398 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 2.480 1.235 3.285 ;
        RECT  0.420 2.480 1.005 2.710 ;
        RECT  0.140 1.210 0.420 2.710 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 3.685 2.240 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.235 1.715 1.570 2.055 ;
        RECT  1.005 0.640 1.235 2.055 ;
        RECT  0.670 1.715 1.005 2.055 ;
    END
END GTIEHBWP7T

MACRO GTIELBWP7T
    CLASS CORE ;
    FOREIGN GTIELBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 0.5400 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 0.640 1.235 1.440 ;
        RECT  0.420 1.210 1.005 1.440 ;
        RECT  0.140 1.210 0.420 2.710 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 3.685 2.240 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.235 1.715 1.570 2.055 ;
        RECT  1.005 1.715 1.235 3.280 ;
        RECT  0.670 1.715 1.005 2.055 ;
    END
END GTIELBWP7T

MACRO GXNR2D1BWP7T
    CLASS CORE ;
    FOREIGN GXNR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 0.695 0.520 0.925 ;
        RECT  0.420 2.995 0.520 3.225 ;
        RECT  0.140 0.695 0.420 3.225 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  1.185 1.820 2.150 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  2.850 1.820 6.160 2.100 ;
        LAYER METAL1 ;
        RECT  5.810 1.715 6.090 2.710 ;
        RECT  5.180 2.330 5.810 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 -0.235 6.720 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  1.310 -0.235 5.410 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 3.685 6.720 4.155 ;
        RECT  5.410 2.995 5.790 4.155 ;
        RECT  1.310 3.685 5.410 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.320 0.640 6.550 3.225 ;
        RECT  6.255 0.640 6.320 1.385 ;
        RECT  6.200 2.995 6.320 3.225 ;
        RECT  3.810 1.155 6.255 1.385 ;
        RECT  4.335 1.770 5.435 2.000 ;
        RECT  4.610 2.905 5.050 3.420 ;
        RECT  3.960 0.695 5.000 0.925 ;
        RECT  4.055 1.770 4.335 3.225 ;
        RECT  3.945 2.940 4.055 3.225 ;
        RECT  3.580 1.155 3.810 2.055 ;
        RECT  3.240 0.695 3.530 0.925 ;
        RECT  3.245 2.380 3.475 3.280 ;
        RECT  2.845 1.615 3.315 2.150 ;
        RECT  2.615 2.380 3.245 2.660 ;
        RECT  3.010 0.695 3.240 1.385 ;
        RECT  2.615 1.155 3.010 1.385 ;
        RECT  2.375 2.905 2.815 3.420 ;
        RECT  2.080 0.695 2.760 0.925 ;
        RECT  2.335 1.155 2.615 2.660 ;
        RECT  1.800 0.695 2.080 3.225 ;
        RECT  1.720 0.695 1.800 0.925 ;
        RECT  1.650 2.940 1.800 3.225 ;
        RECT  1.260 1.535 1.570 2.300 ;
        RECT  0.670 1.210 0.950 2.145 ;
        LAYER VIA12 ;
        RECT  5.820 1.830 6.080 2.090 ;
        RECT  4.690 2.950 4.950 3.210 ;
        RECT  4.065 2.390 4.325 2.650 ;
        RECT  2.910 1.830 3.170 2.090 ;
        RECT  2.460 2.950 2.720 3.210 ;
        RECT  2.345 1.270 2.605 1.530 ;
        RECT  1.810 2.390 2.070 2.650 ;
        RECT  1.280 1.830 1.540 2.090 ;
        RECT  0.680 1.270 0.940 1.530 ;
        LAYER METAL2 ;
        RECT  2.400 2.940 5.010 3.220 ;
        RECT  1.750 2.380 4.385 2.660 ;
        RECT  0.620 1.260 2.670 1.540 ;
    END
END GXNR2D1BWP7T

MACRO GXNR2D2BWP7T
    CLASS CORE ;
    FOREIGN GXNR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 0.640 1.235 1.440 ;
        RECT  1.005 2.480 1.235 3.280 ;
        RECT  0.420 1.210 1.005 1.440 ;
        RECT  0.420 2.480 1.005 2.710 ;
        RECT  0.140 1.210 0.420 2.710 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  2.860 1.820 3.895 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  5.090 1.820 8.400 2.100 ;
        LAYER METAL1 ;
        RECT  8.050 1.715 8.330 2.710 ;
        RECT  7.420 2.330 8.050 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 -0.235 8.960 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  3.550 -0.235 7.650 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.080 -0.235 3.170 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 3.685 8.960 4.155 ;
        RECT  7.650 2.995 8.030 4.155 ;
        RECT  3.550 3.685 7.650 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.560 0.640 8.790 3.225 ;
        RECT  8.495 0.640 8.560 1.385 ;
        RECT  8.440 2.995 8.560 3.225 ;
        RECT  6.050 1.155 8.495 1.385 ;
        RECT  6.575 1.770 7.675 2.000 ;
        RECT  6.840 2.915 7.300 3.415 ;
        RECT  6.200 0.695 7.240 0.925 ;
        RECT  6.295 1.770 6.575 3.225 ;
        RECT  6.185 2.940 6.295 3.225 ;
        RECT  5.820 1.155 6.050 2.100 ;
        RECT  5.480 0.695 5.770 0.925 ;
        RECT  5.485 2.380 5.715 3.280 ;
        RECT  5.085 1.615 5.555 2.150 ;
        RECT  4.855 2.380 5.485 2.660 ;
        RECT  5.250 0.695 5.480 1.385 ;
        RECT  4.855 1.155 5.250 1.385 ;
        RECT  4.620 2.915 5.080 3.415 ;
        RECT  4.345 0.640 5.000 0.925 ;
        RECT  4.575 1.155 4.855 2.660 ;
        RECT  4.065 0.640 4.345 3.225 ;
        RECT  4.015 0.640 4.065 1.385 ;
        RECT  3.910 2.940 4.065 3.225 ;
        RECT  2.705 1.155 4.015 1.385 ;
        RECT  2.910 1.715 3.810 2.150 ;
        RECT  2.400 2.370 2.835 3.275 ;
        RECT  2.475 0.640 2.705 1.385 ;
        RECT  1.700 1.210 2.080 2.055 ;
        RECT  0.670 1.715 1.700 2.055 ;
        LAYER VIA12 ;
        RECT  8.060 1.830 8.320 2.090 ;
        RECT  6.935 2.950 7.195 3.210 ;
        RECT  6.305 2.390 6.565 2.650 ;
        RECT  5.150 1.830 5.410 2.090 ;
        RECT  4.700 2.950 4.960 3.210 ;
        RECT  4.585 1.270 4.845 1.530 ;
        RECT  4.075 2.390 4.335 2.650 ;
        RECT  3.215 1.830 3.475 2.090 ;
        RECT  2.485 2.390 2.745 2.650 ;
        RECT  1.760 1.270 2.020 1.530 ;
        LAYER METAL2 ;
        RECT  4.640 2.940 7.265 3.220 ;
        RECT  2.400 2.380 6.625 2.660 ;
        RECT  1.700 1.260 4.905 1.540 ;
    END
END GXNR2D2BWP7T

MACRO GXOR2D1BWP7T
    CLASS CORE ;
    FOREIGN GXOR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2561 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 0.695 0.520 0.925 ;
        RECT  0.420 2.995 0.520 3.225 ;
        RECT  0.140 0.695 0.420 3.225 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  1.130 1.820 2.150 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.260 6.050 2.055 ;
        RECT  3.810 1.260 5.740 1.540 ;
        RECT  3.580 1.260 3.810 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 -0.235 6.720 0.235 ;
        RECT  5.410 -0.235 5.790 0.925 ;
        RECT  1.310 -0.235 5.410 0.235 ;
        RECT  0.930 -0.235 1.310 0.925 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.790 3.685 6.720 4.155 ;
        RECT  5.410 2.995 5.790 4.155 ;
        RECT  1.310 3.685 5.410 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.300 0.695 6.580 3.225 ;
        RECT  6.200 0.695 6.300 0.925 ;
        RECT  6.200 2.995 6.300 3.225 ;
        RECT  4.335 1.770 5.435 2.000 ;
        RECT  4.620 2.890 5.040 3.420 ;
        RECT  3.960 0.695 5.000 0.925 ;
        RECT  4.055 1.770 4.335 3.225 ;
        RECT  3.945 2.940 4.055 3.225 ;
        RECT  3.240 0.695 3.530 0.925 ;
        RECT  3.245 2.380 3.475 3.280 ;
        RECT  2.845 1.615 3.315 2.150 ;
        RECT  2.615 2.380 3.245 2.660 ;
        RECT  3.010 0.695 3.240 1.385 ;
        RECT  2.615 1.155 3.010 1.385 ;
        RECT  2.390 2.890 2.810 3.420 ;
        RECT  2.080 0.695 2.760 0.925 ;
        RECT  2.335 1.155 2.615 2.660 ;
        RECT  1.800 0.695 2.080 3.225 ;
        RECT  1.720 0.695 1.800 0.925 ;
        RECT  1.650 2.940 1.800 3.225 ;
        RECT  1.260 1.465 1.570 2.205 ;
        RECT  0.670 1.205 0.950 2.120 ;
        LAYER VIA12 ;
        RECT  6.310 1.880 6.570 2.140 ;
        RECT  4.700 2.950 4.960 3.210 ;
        RECT  4.065 2.390 4.325 2.650 ;
        RECT  2.910 1.830 3.170 2.090 ;
        RECT  2.465 2.950 2.725 3.210 ;
        RECT  2.345 1.270 2.605 1.530 ;
        RECT  1.810 2.390 2.070 2.650 ;
        RECT  1.285 1.830 1.545 2.090 ;
        RECT  0.680 1.270 0.940 1.530 ;
        LAYER METAL2 ;
        RECT  6.300 1.820 6.580 2.200 ;
        RECT  2.850 1.820 6.300 2.100 ;
        RECT  2.390 2.940 5.020 3.220 ;
        RECT  1.750 2.380 4.385 2.660 ;
        RECT  0.620 1.260 2.665 1.540 ;
    END
END GXOR2D1BWP7T

MACRO GXOR2D2BWP7T
    CLASS CORE ;
    FOREIGN GXOR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE gacore7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 0.640 1.235 1.440 ;
        RECT  1.005 2.480 1.235 3.280 ;
        RECT  0.420 1.210 1.005 1.440 ;
        RECT  0.420 2.480 1.005 2.710 ;
        RECT  0.140 1.210 0.420 2.710 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL2 ;
        RECT  2.825 1.820 3.880 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.260 8.290 2.055 ;
        RECT  6.050 1.260 7.980 1.540 ;
        RECT  5.820 1.260 6.050 2.055 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 -0.235 8.960 0.235 ;
        RECT  7.650 -0.235 8.030 0.925 ;
        RECT  3.550 -0.235 7.650 0.235 ;
        RECT  3.170 -0.235 3.550 0.925 ;
        RECT  2.080 -0.235 3.170 0.235 ;
        RECT  1.700 -0.235 2.080 0.925 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.925 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 3.685 8.960 4.155 ;
        RECT  7.650 2.995 8.030 4.155 ;
        RECT  3.550 3.685 7.650 4.155 ;
        RECT  3.170 2.995 3.550 4.155 ;
        RECT  2.080 3.685 3.170 4.155 ;
        RECT  1.700 2.995 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.995 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.540 0.695 8.820 3.225 ;
        RECT  8.440 0.695 8.540 0.925 ;
        RECT  8.440 2.995 8.540 3.225 ;
        RECT  6.575 1.770 7.675 2.000 ;
        RECT  6.840 2.790 7.315 3.380 ;
        RECT  6.200 0.695 7.240 0.925 ;
        RECT  6.295 1.770 6.575 3.225 ;
        RECT  6.185 2.940 6.295 3.225 ;
        RECT  5.480 0.695 5.770 0.925 ;
        RECT  5.485 2.380 5.715 3.280 ;
        RECT  5.085 1.615 5.555 2.150 ;
        RECT  4.855 2.380 5.485 2.660 ;
        RECT  5.250 0.695 5.480 1.385 ;
        RECT  4.855 1.155 5.250 1.385 ;
        RECT  4.600 2.890 5.040 3.430 ;
        RECT  4.300 0.640 5.000 0.925 ;
        RECT  4.575 1.155 4.855 2.660 ;
        RECT  4.065 0.640 4.300 3.225 ;
        RECT  4.015 0.640 4.065 1.390 ;
        RECT  2.705 2.380 4.065 2.660 ;
        RECT  3.910 2.940 4.065 3.225 ;
        RECT  2.705 1.160 4.015 1.390 ;
        RECT  2.910 1.715 3.810 2.140 ;
        RECT  2.475 0.640 2.705 1.390 ;
        RECT  2.475 2.380 2.705 3.330 ;
        RECT  1.670 1.210 1.950 2.055 ;
        RECT  0.670 1.715 1.670 2.055 ;
        LAYER VIA12 ;
        RECT  8.550 1.880 8.810 2.140 ;
        RECT  6.935 2.950 7.195 3.210 ;
        RECT  6.305 2.390 6.565 2.650 ;
        RECT  5.225 1.830 5.485 2.090 ;
        RECT  4.720 2.950 4.980 3.210 ;
        RECT  4.585 1.270 4.845 1.530 ;
        RECT  4.030 2.390 4.290 2.650 ;
        RECT  3.190 1.830 3.450 2.090 ;
        RECT  1.680 1.270 1.940 1.530 ;
        LAYER METAL2 ;
        RECT  8.540 1.820 8.820 2.200 ;
        RECT  5.140 1.820 8.540 2.100 ;
        RECT  4.660 2.940 7.255 3.220 ;
        RECT  3.935 2.380 6.625 2.660 ;
        RECT  1.605 1.260 4.905 1.540 ;
    END
END GXOR2D2BWP7T

MACRO HA1D0BWP7T
    CLASS CORE ;
    FOREIGN HA1D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN S
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.935 0.835 8.260 2.780 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 0.5813 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 0.945 0.465 1.285 ;
        RECT  0.420 2.560 0.465 2.900 ;
        RECT  0.140 0.945 0.420 2.900 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.7371 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.605 3.225 7.005 3.455 ;
        RECT  4.325 2.790 4.605 3.455 ;
        RECT  2.305 2.790 4.325 3.020 ;
        RECT  2.075 1.740 2.305 3.020 ;
        RECT  1.260 1.740 2.075 2.150 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.605 3.830 2.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.445 -0.235 8.400 0.235 ;
        RECT  7.215 -0.235 7.445 1.170 ;
        RECT  3.890 -0.235 7.215 0.235 ;
        RECT  3.510 -0.235 3.890 0.670 ;
        RECT  0.520 -0.235 3.510 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.605 3.685 8.400 4.155 ;
        RECT  7.265 3.455 7.605 4.155 ;
        RECT  3.915 3.685 7.265 4.155 ;
        RECT  3.455 3.250 3.915 4.155 ;
        RECT  2.435 3.685 3.455 4.155 ;
        RECT  2.095 3.455 2.435 4.155 ;
        RECT  1.025 3.685 2.095 4.155 ;
        RECT  0.685 3.455 1.025 4.155 ;
        RECT  0.000 3.685 0.685 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.415 1.600 7.645 2.995 ;
        RECT  5.440 2.765 7.415 2.995 ;
        RECT  6.630 0.890 6.780 1.120 ;
        RECT  6.630 2.300 6.780 2.535 ;
        RECT  6.400 0.890 6.630 2.535 ;
        RECT  6.300 1.685 6.400 2.110 ;
        RECT  5.970 2.300 6.080 2.535 ;
        RECT  5.970 0.925 6.025 1.265 ;
        RECT  5.740 0.465 5.970 2.535 ;
        RECT  4.350 0.465 5.740 0.695 ;
        RECT  5.190 0.925 5.440 2.995 ;
        RECT  5.020 0.925 5.190 1.155 ;
        RECT  4.980 2.760 5.190 2.995 ;
        RECT  4.120 0.465 4.350 2.560 ;
        RECT  2.800 0.900 4.120 1.130 ;
        RECT  2.715 2.330 4.120 2.560 ;
        RECT  0.935 0.695 2.440 0.925 ;
        RECT  0.935 2.680 1.845 2.910 ;
        RECT  0.705 0.695 0.935 2.910 ;
        RECT  0.650 1.790 0.705 2.130 ;
    END
END HA1D0BWP7T

MACRO HA1D1BWP7T
    CLASS CORE ;
    FOREIGN HA1D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN S
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.495 0.930 8.820 2.780 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.365 0.495 0.465 1.305 ;
        RECT  0.365 2.245 0.465 3.350 ;
        RECT  0.135 0.495 0.365 3.350 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.9171 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.235 3.225 7.275 3.455 ;
        RECT  4.955 2.790 5.235 3.455 ;
        RECT  2.440 2.790 4.955 3.020 ;
        RECT  2.210 1.770 2.440 3.020 ;
        RECT  1.210 1.770 2.210 2.150 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 1.2636 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.545 3.830 2.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.005 -0.235 8.960 0.235 ;
        RECT  7.775 -0.235 8.005 1.265 ;
        RECT  4.520 -0.235 7.775 0.235 ;
        RECT  4.140 -0.235 4.520 0.670 ;
        RECT  3.060 -0.235 4.140 0.235 ;
        RECT  2.300 -0.235 3.060 0.465 ;
        RECT  1.265 -0.235 2.300 0.235 ;
        RECT  0.885 -0.235 1.265 0.785 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.965 3.685 8.960 4.155 ;
        RECT  7.625 3.455 7.965 4.155 ;
        RECT  4.545 3.685 7.625 4.155 ;
        RECT  4.085 3.250 4.545 4.155 ;
        RECT  2.720 3.685 4.085 4.155 ;
        RECT  2.380 3.250 2.720 4.155 ;
        RECT  1.255 3.685 2.380 4.155 ;
        RECT  0.875 3.155 1.255 4.155 ;
        RECT  0.000 3.685 0.875 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.975 1.600 8.205 2.995 ;
        RECT  6.000 2.765 7.975 2.995 ;
        RECT  7.190 0.985 7.340 1.215 ;
        RECT  7.190 2.300 7.340 2.535 ;
        RECT  6.960 0.985 7.190 2.535 ;
        RECT  6.860 1.685 6.960 2.110 ;
        RECT  6.530 2.300 6.640 2.535 ;
        RECT  6.530 0.925 6.585 1.265 ;
        RECT  6.300 0.465 6.530 2.535 ;
        RECT  4.980 0.465 6.300 0.695 ;
        RECT  5.750 0.925 6.000 2.995 ;
        RECT  5.580 0.925 5.750 1.155 ;
        RECT  5.540 2.760 5.750 2.995 ;
        RECT  4.750 0.465 4.980 1.130 ;
        RECT  4.675 0.900 4.750 1.130 ;
        RECT  4.445 0.900 4.675 2.560 ;
        RECT  3.430 0.900 4.445 1.130 ;
        RECT  3.430 2.330 4.445 2.560 ;
        RECT  0.925 1.020 2.500 1.250 ;
        RECT  1.675 2.405 1.905 3.220 ;
        RECT  0.925 2.405 1.675 2.635 ;
        RECT  0.695 1.020 0.925 2.635 ;
        RECT  0.595 1.540 0.695 1.880 ;
    END
END HA1D1BWP7T

MACRO HA1D2BWP7T
    CLASS CORE ;
    FOREIGN HA1D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN S
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.740 1.060 9.940 2.490 ;
        RECT  9.660 0.495 9.740 3.315 ;
        RECT  9.455 0.495 9.660 1.345 ;
        RECT  9.455 2.205 9.660 3.315 ;
        END
    END S
    PIN CO
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 0.495 1.185 1.305 ;
        RECT  0.980 2.245 1.185 3.350 ;
        RECT  0.955 0.495 0.980 3.350 ;
        RECT  0.700 0.985 0.955 2.475 ;
        END
    END CO
    PIN B
        ANTENNAGATEAREA 0.9171 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.115 3.225 8.450 3.455 ;
        RECT  5.835 2.790 6.115 3.455 ;
        RECT  3.220 2.790 5.835 3.020 ;
        RECT  2.990 1.770 3.220 3.020 ;
        RECT  1.930 1.770 2.990 2.150 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 1.2636 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 1.545 4.390 2.100 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 -0.235 10.640 0.235 ;
        RECT  10.175 -0.235 10.405 1.305 ;
        RECT  8.945 -0.235 10.175 0.235 ;
        RECT  8.715 -0.235 8.945 0.905 ;
        RECT  5.400 -0.235 8.715 0.235 ;
        RECT  5.020 -0.235 5.400 0.670 ;
        RECT  3.930 -0.235 5.020 0.235 ;
        RECT  3.590 -0.235 3.930 1.140 ;
        RECT  1.985 -0.235 3.590 0.235 ;
        RECT  1.605 -0.235 1.985 0.785 ;
        RECT  0.465 -0.235 1.605 0.235 ;
        RECT  0.235 -0.235 0.465 1.305 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 3.685 10.640 4.155 ;
        RECT  10.175 2.255 10.405 4.155 ;
        RECT  9.020 3.685 10.175 4.155 ;
        RECT  8.680 3.250 9.020 4.155 ;
        RECT  5.425 3.685 8.680 4.155 ;
        RECT  4.965 3.250 5.425 4.155 ;
        RECT  3.440 3.685 4.965 4.155 ;
        RECT  3.100 3.250 3.440 4.155 ;
        RECT  1.975 3.685 3.100 4.155 ;
        RECT  1.595 3.155 1.975 4.155 ;
        RECT  0.465 3.685 1.595 4.155 ;
        RECT  0.235 2.255 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.935 1.600 9.165 2.995 ;
        RECT  6.880 2.765 8.935 2.995 ;
        RECT  8.110 0.585 8.260 0.815 ;
        RECT  8.110 2.300 8.260 2.535 ;
        RECT  7.880 0.585 8.110 2.535 ;
        RECT  7.780 1.685 7.880 2.110 ;
        RECT  7.410 2.300 7.520 2.535 ;
        RECT  7.410 0.925 7.465 1.265 ;
        RECT  7.180 0.465 7.410 2.535 ;
        RECT  5.860 0.465 7.180 0.695 ;
        RECT  6.630 0.925 6.880 2.995 ;
        RECT  6.460 0.925 6.630 1.155 ;
        RECT  6.420 2.760 6.630 2.995 ;
        RECT  5.630 0.465 5.860 1.130 ;
        RECT  5.555 0.900 5.630 1.130 ;
        RECT  5.325 0.900 5.555 2.560 ;
        RECT  4.310 0.900 5.325 1.130 ;
        RECT  4.040 2.330 5.325 2.560 ;
        RECT  1.645 1.020 3.220 1.250 ;
        RECT  2.395 2.405 2.625 3.220 ;
        RECT  1.645 2.405 2.395 2.635 ;
        RECT  1.415 1.020 1.645 2.635 ;
        RECT  1.315 1.540 1.415 1.880 ;
    END
END HA1D2BWP7T

MACRO IAO21D0BWP7T
    CLASS CORE ;
    FOREIGN IAO21D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6296 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.825 3.220 3.285 ;
        RECT  2.180 0.825 2.940 1.055 ;
        RECT  2.840 3.055 2.940 3.285 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 2.700 2.710 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 1.770 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.455 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.815 -0.235 3.360 0.235 ;
        RECT  1.435 -0.235 1.815 1.055 ;
        RECT  0.000 -0.235 1.435 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.870 3.685 3.360 4.155 ;
        RECT  1.490 3.030 1.870 4.155 ;
        RECT  0.000 3.685 1.490 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.910 1.300 2.140 1.920 ;
        RECT  1.030 1.300 1.910 1.540 ;
        RECT  0.945 0.770 1.030 1.540 ;
        RECT  0.705 0.770 0.945 3.185 ;
        RECT  0.180 2.955 0.705 3.185 ;
    END
END IAO21D0BWP7T

MACRO IAO21D1BWP7T
    CLASS CORE ;
    FOREIGN IAO21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.120 3.780 2.710 ;
        RECT  2.795 1.120 3.500 1.360 ;
        RECT  3.395 2.310 3.500 2.710 ;
        RECT  3.165 2.310 3.395 3.425 ;
        RECT  2.565 0.670 2.795 1.360 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.765 1.735 3.040 1.970 ;
        RECT  2.480 1.735 2.765 2.710 ;
        RECT  1.820 2.330 2.480 2.710 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2484 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.730 1.545 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2484 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.630 -0.235 3.920 0.235 ;
        RECT  3.250 -0.235 3.630 0.880 ;
        RECT  2.090 -0.235 3.250 0.235 ;
        RECT  1.710 -0.235 2.090 0.770 ;
        RECT  0.650 -0.235 1.710 0.235 ;
        RECT  0.270 -0.235 0.650 0.740 ;
        RECT  0.000 -0.235 0.270 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.010 3.685 3.920 4.155 ;
        RECT  1.630 3.060 2.010 4.155 ;
        RECT  0.000 3.685 1.630 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.975 1.220 2.205 2.000 ;
        RECT  1.295 1.220 1.975 1.460 ;
        RECT  1.065 0.525 1.295 1.460 ;
        RECT  0.965 1.220 1.065 1.460 ;
        RECT  0.725 1.220 0.965 3.305 ;
        RECT  0.290 3.075 0.725 3.305 ;
    END
END IAO21D1BWP7T

MACRO IAO21D2BWP7T
    CLASS CORE ;
    FOREIGN IAO21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8198 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.840 0.495 4.070 1.370 ;
        RECT  3.780 1.120 3.840 1.370 ;
        RECT  3.500 1.120 3.780 2.755 ;
        RECT  2.630 1.120 3.500 1.400 ;
        RECT  3.065 2.520 3.500 2.755 ;
        RECT  2.400 0.495 2.630 1.400 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.670 3.220 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.600 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.170 0.450 2.190 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.865 -0.235 5.040 0.235 ;
        RECT  4.485 -0.235 4.865 1.200 ;
        RECT  3.430 -0.235 4.485 0.235 ;
        RECT  3.050 -0.235 3.430 0.880 ;
        RECT  1.985 -0.235 3.050 0.235 ;
        RECT  1.605 -0.235 1.985 0.785 ;
        RECT  0.540 -0.235 1.605 0.235 ;
        RECT  0.160 -0.235 0.540 0.785 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.790 3.685 5.040 4.155 ;
        RECT  4.560 2.245 4.790 4.155 ;
        RECT  1.905 3.685 4.560 4.155 ;
        RECT  1.525 3.065 1.905 4.155 ;
        RECT  0.000 3.685 1.525 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.055 1.650 4.285 3.270 ;
        RECT  2.650 3.030 4.055 3.270 ;
        RECT  2.410 2.505 2.650 3.270 ;
        RECT  2.130 2.505 2.410 2.745 ;
        RECT  1.900 1.100 2.130 2.745 ;
        RECT  1.195 1.100 1.900 1.340 ;
        RECT  0.955 0.465 1.195 1.340 ;
        RECT  0.935 1.100 0.955 1.340 ;
        RECT  0.690 1.100 0.935 2.700 ;
        RECT  0.475 2.470 0.690 2.700 ;
        RECT  0.230 2.470 0.475 3.380 ;
    END
END IAO21D2BWP7T

MACRO IAO22D0BWP7T
    CLASS CORE ;
    FOREIGN IAO22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.7792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 0.640 4.245 1.240 ;
        RECT  2.660 0.640 4.015 0.880 ;
        RECT  2.385 0.640 2.660 2.905 ;
        RECT  2.380 0.955 2.385 2.905 ;
        RECT  2.005 0.955 2.380 1.185 ;
        RECT  2.005 2.675 2.380 2.905 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.245 2.190 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 4.345 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.080 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.850 -0.235 4.480 0.235 ;
        RECT  1.485 -0.235 1.850 0.465 ;
        RECT  0.000 -0.235 1.485 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 3.685 4.480 4.155 ;
        RECT  3.365 2.680 3.745 4.155 ;
        RECT  1.835 3.685 3.365 4.155 ;
        RECT  1.475 3.450 1.835 4.155 ;
        RECT  0.000 3.685 1.475 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.605 1.645 2.135 1.985 ;
        RECT  1.365 0.895 1.605 3.190 ;
        RECT  0.745 0.895 1.365 1.125 ;
        RECT  0.465 2.960 1.365 3.190 ;
        RECT  0.235 2.960 0.465 3.430 ;
    END
END IAO22D0BWP7T

MACRO IAO22D1BWP7T
    CLASS CORE ;
    FOREIGN IAO22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.4324 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.625 3.220 2.400 ;
        RECT  2.645 2.160 2.940 2.400 ;
        RECT  2.415 2.160 2.645 3.390 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.690 4.900 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.730 1.540 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.815 -0.235 5.040 0.235 ;
        RECT  4.565 -0.235 4.815 1.275 ;
        RECT  2.290 -0.235 4.565 0.235 ;
        RECT  1.910 -0.235 2.290 0.995 ;
        RECT  0.580 -0.235 1.910 0.235 ;
        RECT  0.200 -0.235 0.580 1.095 ;
        RECT  0.000 -0.235 0.200 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.155 3.685 5.040 4.155 ;
        RECT  3.775 3.115 4.155 4.155 ;
        RECT  0.580 3.685 3.775 4.155 ;
        RECT  0.200 2.960 0.580 4.155 ;
        RECT  0.000 3.685 0.200 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.575 2.640 4.805 3.450 ;
        RECT  3.365 2.640 4.575 2.870 ;
        RECT  3.135 2.640 3.365 3.450 ;
        RECT  2.055 1.675 2.630 1.905 ;
        RECT  1.825 1.260 2.055 3.220 ;
        RECT  1.250 1.260 1.825 1.490 ;
        RECT  1.545 2.990 1.825 3.220 ;
        RECT  1.020 0.805 1.250 1.490 ;
    END
END IAO22D1BWP7T

MACRO IAO22D2BWP7T
    CLASS CORE ;
    FOREIGN IAO22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.7250 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.055 4.340 2.710 ;
        RECT  4.055 1.055 4.060 1.295 ;
        RECT  3.455 2.330 4.060 2.710 ;
        RECT  3.825 0.465 4.055 1.295 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.710 1.770 6.020 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.210 4.900 2.530 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.550 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.735 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.845 -0.235 6.160 0.235 ;
        RECT  4.465 -0.235 4.845 0.735 ;
        RECT  3.350 -0.235 4.465 0.235 ;
        RECT  3.010 -0.235 3.350 0.465 ;
        RECT  2.010 -0.235 3.010 0.235 ;
        RECT  1.645 -0.235 2.010 0.465 ;
        RECT  0.000 -0.235 1.645 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 3.685 6.160 4.155 ;
        RECT  5.695 3.040 5.925 4.155 ;
        RECT  4.500 3.685 5.695 4.155 ;
        RECT  4.160 3.455 4.500 4.155 ;
        RECT  2.625 3.685 4.160 4.155 ;
        RECT  2.285 3.455 2.625 4.155 ;
        RECT  0.520 3.685 2.285 4.155 ;
        RECT  0.180 3.455 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.465 0.480 5.980 0.710 ;
        RECT  5.235 0.480 5.465 3.210 ;
        RECT  0.570 2.980 5.235 3.210 ;
        RECT  3.175 1.725 3.780 1.955 ;
        RECT  2.945 1.725 3.175 2.745 ;
        RECT  1.030 2.515 2.945 2.745 ;
        RECT  2.420 0.695 2.760 1.115 ;
        RECT  1.185 0.695 2.420 0.925 ;
        RECT  0.955 0.485 1.185 0.925 ;
        RECT  0.800 1.155 1.030 2.745 ;
        RECT  0.465 1.155 0.800 1.385 ;
        RECT  0.340 1.670 0.570 3.210 ;
        RECT  0.235 0.465 0.465 1.385 ;
    END
END IAO22D2BWP7T

MACRO IIND4D0BWP7T
    CLASS CORE ;
    FOREIGN IIND4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.135 2.725 3.365 3.370 ;
        RECT  2.100 2.725 3.135 2.955 ;
        RECT  1.910 0.880 2.100 2.955 ;
        RECT  1.820 0.880 1.910 3.350 ;
        RECT  1.555 0.880 1.820 1.220 ;
        RECT  1.680 2.725 1.820 3.350 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.495 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.650 2.695 1.820 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 1.210 4.900 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.585 -0.235 5.040 0.235 ;
        RECT  1.220 -0.235 1.585 0.465 ;
        RECT  0.000 -0.235 1.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.165 3.685 5.040 4.155 ;
        RECT  3.785 2.920 4.165 4.155 ;
        RECT  2.715 3.685 3.785 4.155 ;
        RECT  2.335 3.185 2.715 4.155 ;
        RECT  1.280 3.685 2.335 4.155 ;
        RECT  0.900 2.915 1.280 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.325 0.700 4.860 0.930 ;
        RECT  4.575 2.380 4.805 3.205 ;
        RECT  4.325 2.380 4.575 2.610 ;
        RECT  4.085 0.700 4.325 2.610 ;
        RECT  3.630 1.760 4.085 2.100 ;
        RECT  1.005 0.725 1.235 2.630 ;
        RECT  0.465 0.725 1.005 0.955 ;
        RECT  0.470 2.390 1.005 2.630 ;
        RECT  0.235 2.390 0.470 3.205 ;
        RECT  0.235 0.500 0.465 0.955 ;
    END
END IIND4D0BWP7T

MACRO IIND4D1BWP7T
    CLASS CORE ;
    FOREIGN IIND4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.9596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 2.475 3.730 3.325 ;
        RECT  2.100 2.475 3.500 2.715 ;
        RECT  1.905 0.590 2.100 2.715 ;
        RECT  1.820 0.590 1.905 3.335 ;
        RECT  1.615 0.590 1.820 0.825 ;
        RECT  1.675 2.420 1.820 3.335 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        RECT  3.205 1.695 3.500 1.925 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.670 1.595 2.875 1.825 ;
        RECT  2.380 0.650 2.670 1.825 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.210 5.460 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.190 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 -0.235 5.600 0.235 ;
        RECT  4.220 -0.235 4.450 0.785 ;
        RECT  0.540 -0.235 4.220 0.235 ;
        RECT  0.160 -0.235 0.540 0.710 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 3.685 5.600 4.155 ;
        RECT  4.240 3.060 4.620 4.155 ;
        RECT  2.865 3.685 4.240 4.155 ;
        RECT  2.485 2.990 2.865 4.155 ;
        RECT  1.260 3.685 2.485 4.155 ;
        RECT  0.880 3.055 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.920 0.480 5.420 0.710 ;
        RECT  5.135 2.545 5.365 3.380 ;
        RECT  4.920 2.545 5.135 2.775 ;
        RECT  4.690 0.480 4.920 2.775 ;
        RECT  4.040 1.685 4.690 1.915 ;
        RECT  0.955 0.465 1.200 2.745 ;
        RECT  0.465 2.505 0.955 2.745 ;
        RECT  0.235 2.505 0.465 3.395 ;
    END
END IIND4D1BWP7T

MACRO IIND4D2BWP7T
    CLASS CORE ;
    FOREIGN IIND4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.4992 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 2.515 8.460 2.745 ;
        RECT  3.500 0.955 3.780 2.745 ;
        RECT  3.120 0.955 3.500 1.185 ;
        RECT  3.225 2.515 3.500 2.745 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.625 7.140 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.625 5.460 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.600 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.580 -0.235 9.520 0.235 ;
        RECT  8.200 -0.235 8.580 0.840 ;
        RECT  1.305 -0.235 8.200 0.235 ;
        RECT  0.925 -0.235 1.305 0.825 ;
        RECT  0.000 -0.235 0.925 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.240 3.685 9.520 4.155 ;
        RECT  8.870 3.455 9.240 4.155 ;
        RECT  7.645 3.685 8.870 4.155 ;
        RECT  7.285 3.455 7.645 4.155 ;
        RECT  6.055 3.685 7.285 4.155 ;
        RECT  5.710 3.455 6.055 4.155 ;
        RECT  4.375 3.685 5.710 4.155 ;
        RECT  4.030 3.455 4.375 4.155 ;
        RECT  2.805 3.685 4.030 4.155 ;
        RECT  2.460 3.455 2.805 4.155 ;
        RECT  1.280 3.685 2.460 4.155 ;
        RECT  0.930 3.455 1.280 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.995 0.495 9.225 1.360 ;
        RECT  8.890 1.700 9.120 3.220 ;
        RECT  7.790 1.110 8.995 1.360 ;
        RECT  7.965 1.700 8.890 1.930 ;
        RECT  1.000 2.980 8.890 3.220 ;
        RECT  7.555 0.465 7.790 1.360 ;
        RECT  6.345 0.465 7.555 0.705 ;
        RECT  6.835 0.965 7.065 1.360 ;
        RECT  4.895 1.120 6.835 1.360 ;
        RECT  6.115 0.465 6.345 0.840 ;
        RECT  5.385 0.465 5.615 0.840 ;
        RECT  2.685 0.465 5.385 0.705 ;
        RECT  4.665 0.965 4.895 1.360 ;
        RECT  2.135 1.665 3.075 1.900 ;
        RECT  2.455 0.465 2.685 1.305 ;
        RECT  1.905 0.635 2.135 2.745 ;
        RECT  1.700 0.635 1.905 0.865 ;
        RECT  1.765 2.515 1.905 2.745 ;
        RECT  0.760 1.090 1.000 3.220 ;
        RECT  0.465 1.090 0.760 1.320 ;
        RECT  0.180 2.980 0.760 3.220 ;
        RECT  0.235 0.495 0.465 1.320 ;
    END
END IIND4D2BWP7T

MACRO IINR4D0BWP7T
    CLASS CORE ;
    FOREIGN IINR4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1008 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.120 0.475 3.350 1.220 ;
        RECT  1.905 0.990 3.120 1.220 ;
        RECT  1.820 2.290 2.100 3.455 ;
        RECT  1.755 0.475 1.905 1.220 ;
        RECT  1.755 2.290 1.820 2.660 ;
        RECT  1.170 3.225 1.820 3.455 ;
        RECT  1.675 0.475 1.755 2.660 ;
        RECT  1.525 0.990 1.675 2.660 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 1.725 3.830 2.065 ;
        RECT  3.500 1.725 3.780 2.750 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.500 3.220 2.750 ;
        RECT  2.825 1.500 2.940 1.730 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 2.385 4.465 2.750 ;
        RECT  4.060 1.770 4.340 2.750 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.475 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.155 -0.235 5.040 0.235 ;
        RECT  3.775 -0.235 4.155 0.760 ;
        RECT  2.685 -0.235 3.775 0.235 ;
        RECT  2.345 -0.235 2.685 0.760 ;
        RECT  1.255 -0.235 2.345 0.235 ;
        RECT  0.875 -0.235 1.255 0.760 ;
        RECT  0.000 -0.235 0.875 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.115 3.685 5.040 4.155 ;
        RECT  3.735 3.455 4.115 4.155 ;
        RECT  0.725 3.685 3.735 4.155 ;
        RECT  0.385 3.455 0.725 4.155 ;
        RECT  0.000 3.685 0.385 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.695 0.530 4.925 3.225 ;
        RECT  4.510 0.530 4.695 0.760 ;
        RECT  2.595 2.995 4.695 3.225 ;
        RECT  2.365 1.450 2.595 3.225 ;
        RECT  2.155 1.450 2.365 1.680 ;
        RECT  1.040 1.120 1.270 2.645 ;
        RECT  0.465 1.120 1.040 1.360 ;
        RECT  0.745 2.415 1.040 2.645 ;
        RECT  0.235 0.475 0.465 1.360 ;
    END
END IINR4D0BWP7T

MACRO IINR4D1BWP7T
    CLASS CORE ;
    FOREIGN IINR4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.7538 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 2.380 4.050 2.660 ;
        RECT  3.565 0.595 3.795 0.935 ;
        RECT  2.885 0.695 3.565 0.935 ;
        RECT  2.655 0.695 2.885 2.660 ;
        RECT  1.185 0.695 2.655 0.925 ;
        RECT  0.955 0.585 1.185 0.925 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.425 1.210 1.540 1.590 ;
        RECT  1.195 1.210 1.425 1.825 ;
        RECT  0.700 1.210 1.195 1.590 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.220 2.375 2.340 ;
        RECT  0.465 2.100 2.145 2.340 ;
        RECT  0.140 1.210 0.465 2.340 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 0.700 6.070 0.980 ;
        RECT  5.735 0.700 6.020 1.630 ;
        RECT  5.690 0.700 5.735 0.980 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.170 6.635 2.190 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.315 -0.235 7.280 0.235 ;
        RECT  5.975 -0.235 6.315 0.465 ;
        RECT  4.570 -0.235 5.975 0.235 ;
        RECT  4.230 -0.235 4.570 0.965 ;
        RECT  3.090 -0.235 4.230 0.235 ;
        RECT  2.750 -0.235 3.090 0.465 ;
        RECT  2.000 -0.235 2.750 0.235 ;
        RECT  1.660 -0.235 2.000 0.465 ;
        RECT  0.520 -0.235 1.660 0.235 ;
        RECT  0.180 -0.235 0.520 0.670 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.280 3.685 7.280 4.155 ;
        RECT  5.940 3.455 6.280 4.155 ;
        RECT  1.740 3.685 5.940 4.155 ;
        RECT  1.360 3.140 1.740 4.155 ;
        RECT  0.000 3.685 1.360 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.900 0.570 7.140 2.995 ;
        RECT  6.760 0.570 6.900 0.810 ;
        RECT  6.810 2.460 6.900 2.995 ;
        RECT  4.595 2.765 6.810 2.995 ;
        RECT  5.185 2.305 5.740 2.535 ;
        RECT  5.185 0.575 5.355 0.805 ;
        RECT  2.280 3.225 5.245 3.455 ;
        RECT  4.955 0.575 5.185 2.535 ;
        RECT  3.130 1.240 4.955 1.470 ;
        RECT  3.930 1.780 4.355 2.010 ;
        RECT  2.050 2.635 2.280 3.455 ;
        RECT  0.465 2.635 2.050 2.865 ;
        RECT  0.235 2.635 0.465 3.445 ;
        RECT  4.355 1.780 4.595 2.995 ;
    END
END IINR4D1BWP7T

MACRO IINR4D2BWP7T
    CLASS CORE ;
    FOREIGN IINR4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.6596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.995 0.700 12.760 0.930 ;
        RECT  5.765 0.700 5.995 1.415 ;
        RECT  3.780 1.185 5.765 1.415 ;
        RECT  3.780 2.250 3.890 2.885 ;
        RECT  3.660 1.185 3.780 2.885 ;
        RECT  3.500 1.185 3.660 2.490 ;
        RECT  2.755 1.185 3.500 1.415 ;
        RECT  2.450 2.250 3.500 2.490 ;
        RECT  2.520 0.485 2.755 1.415 ;
        RECT  2.220 2.250 2.450 2.910 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.490 1.690 13.710 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.595 1.690 10.815 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.215 1.690 15.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.475 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.495 -0.235 15.680 0.235 ;
        RECT  15.155 -0.235 15.495 1.195 ;
        RECT  13.540 -0.235 15.155 0.235 ;
        RECT  13.200 -0.235 13.540 0.785 ;
        RECT  11.920 -0.235 13.200 0.235 ;
        RECT  11.580 -0.235 11.920 0.470 ;
        RECT  10.720 -0.235 11.580 0.235 ;
        RECT  10.380 -0.235 10.720 0.470 ;
        RECT  9.030 -0.235 10.380 0.235 ;
        RECT  8.690 -0.235 9.030 0.470 ;
        RECT  6.970 -0.235 8.690 0.235 ;
        RECT  6.630 -0.235 6.970 0.465 ;
        RECT  5.365 -0.235 6.630 0.235 ;
        RECT  4.985 -0.235 5.365 0.920 ;
        RECT  3.585 -0.235 4.985 0.235 ;
        RECT  3.205 -0.235 3.585 0.920 ;
        RECT  2.085 -0.235 3.205 0.235 ;
        RECT  1.745 -0.235 2.085 1.200 ;
        RECT  0.525 -0.235 1.745 0.235 ;
        RECT  0.185 -0.235 0.525 0.825 ;
        RECT  0.000 -0.235 0.185 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.500 3.685 15.680 4.155 ;
        RECT  15.160 3.040 15.500 4.155 ;
        RECT  13.480 3.685 15.160 4.155 ;
        RECT  13.140 2.840 13.480 4.155 ;
        RECT  12.040 3.685 13.140 4.155 ;
        RECT  11.700 2.840 12.040 4.155 ;
        RECT  0.525 3.685 11.700 4.155 ;
        RECT  0.185 2.505 0.525 4.155 ;
        RECT  0.000 3.685 0.185 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.455 0.495 14.685 3.450 ;
        RECT  7.820 1.190 14.455 1.420 ;
        RECT  12.705 2.380 14.200 2.610 ;
        RECT  12.475 2.380 12.705 3.310 ;
        RECT  11.265 2.380 12.475 2.610 ;
        RECT  11.035 2.380 11.265 3.455 ;
        RECT  9.825 3.225 11.035 3.455 ;
        RECT  10.315 2.380 10.550 2.885 ;
        RECT  9.105 2.380 10.315 2.610 ;
        RECT  9.595 2.860 9.825 3.455 ;
        RECT  8.385 3.225 9.595 3.455 ;
        RECT  8.875 2.380 9.105 2.885 ;
        RECT  6.770 2.380 8.875 2.610 ;
        RECT  8.155 2.860 8.385 3.455 ;
        RECT  7.590 1.190 7.820 1.925 ;
        RECT  4.825 1.690 7.590 1.925 ;
        RECT  7.255 2.890 7.490 3.455 ;
        RECT  6.050 3.225 7.255 3.455 ;
        RECT  6.540 2.380 6.770 2.885 ;
        RECT  5.330 2.380 6.540 2.610 ;
        RECT  5.820 2.890 6.050 3.455 ;
        RECT  4.610 3.225 5.820 3.455 ;
        RECT  5.100 2.380 5.330 2.885 ;
        RECT  4.380 2.525 4.610 3.455 ;
        RECT  3.170 3.225 4.380 3.455 ;
        RECT  1.190 1.695 3.220 1.925 ;
        RECT  2.940 2.740 3.170 3.455 ;
        RECT  1.730 3.225 2.940 3.455 ;
        RECT  1.500 3.110 1.730 3.455 ;
        RECT  0.960 0.485 1.190 2.705 ;
    END
END IINR4D2BWP7T

MACRO IND2D0BWP7T
    CLASS CORE ;
    FOREIGN IND2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6099 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.575 2.660 2.710 ;
        RECT  2.205 0.575 2.380 0.805 ;
        RECT  1.505 2.480 2.380 2.710 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.730 0.465 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 -0.235 2.800 0.235 ;
        RECT  0.880 -0.235 1.260 0.765 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.605 3.685 2.800 4.155 ;
        RECT  2.265 2.980 2.605 4.155 ;
        RECT  1.525 3.685 2.265 4.155 ;
        RECT  1.160 3.455 1.525 4.155 ;
        RECT  0.000 3.685 1.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.945 1.655 1.475 1.885 ;
        RECT  0.935 1.170 0.945 1.885 ;
        RECT  0.705 1.170 0.935 3.345 ;
        RECT  0.465 1.170 0.705 1.410 ;
        RECT  0.180 3.115 0.705 3.345 ;
        RECT  0.235 0.480 0.465 1.410 ;
    END
END IND2D0BWP7T

MACRO IND2D1BWP7T
    CLASS CORE ;
    FOREIGN IND2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2198 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 0.655 2.620 0.885 ;
        RECT  1.845 0.655 2.100 2.750 ;
        RECT  1.820 0.655 1.845 3.350 ;
        RECT  1.615 2.360 1.820 3.350 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.210 2.660 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.470 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 -0.235 2.800 0.235 ;
        RECT  0.935 -0.235 1.290 0.465 ;
        RECT  0.000 -0.235 0.935 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.565 3.685 2.800 4.155 ;
        RECT  2.335 2.490 2.565 4.155 ;
        RECT  1.080 3.685 2.335 4.155 ;
        RECT  0.725 3.440 1.080 4.155 ;
        RECT  0.000 3.685 0.725 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.195 1.690 1.540 1.925 ;
        RECT  0.965 0.700 1.195 2.660 ;
        RECT  0.180 0.700 0.965 0.930 ;
        RECT  0.180 2.430 0.965 2.660 ;
    END
END IND2D1BWP7T

MACRO IND2D2BWP7T
    CLASS CORE ;
    FOREIGN IND2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.0196 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.735 4.340 2.850 ;
        RECT  2.340 0.735 4.060 0.965 ;
        RECT  3.345 2.620 4.060 2.850 ;
        RECT  3.115 2.620 3.345 3.430 ;
        RECT  1.910 2.620 3.115 2.850 ;
        RECT  1.675 2.620 1.910 3.430 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.715 2.920 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 -0.235 4.480 0.235 ;
        RECT  3.750 -0.235 4.100 0.465 ;
        RECT  1.285 -0.235 3.750 0.235 ;
        RECT  0.925 -0.235 1.285 0.470 ;
        RECT  0.000 -0.235 0.925 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 3.685 4.480 4.155 ;
        RECT  3.760 3.140 4.140 4.155 ;
        RECT  2.700 3.685 3.760 4.155 ;
        RECT  2.320 3.140 2.700 4.155 ;
        RECT  1.260 3.685 2.320 4.155 ;
        RECT  0.880 2.940 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 1.935 ;
        RECT  1.585 1.210 3.500 1.450 ;
        RECT  1.355 1.210 1.585 1.920 ;
        RECT  0.990 1.690 1.355 1.920 ;
        RECT  0.760 0.750 0.990 2.680 ;
        RECT  0.465 0.750 0.760 0.980 ;
        RECT  0.465 2.450 0.760 2.680 ;
        RECT  0.235 0.640 0.465 0.980 ;
        RECT  0.235 2.450 0.465 3.370 ;
    END
END IND2D2BWP7T

MACRO IND2D4BWP7T
    CLASS CORE ;
    FOREIGN IND2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 4.2588 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.155 1.450 7.450 3.105 ;
        RECT  6.970 1.450 7.155 2.835 ;
        RECT  6.550 1.020 6.970 2.835 ;
        RECT  6.310 1.020 6.550 1.250 ;
        RECT  5.840 2.605 6.550 2.835 ;
        RECT  5.600 2.605 5.840 3.415 ;
        RECT  4.225 2.605 5.600 2.835 ;
        RECT  3.995 2.605 4.225 3.405 ;
        RECT  3.140 2.605 3.995 2.835 ;
        RECT  3.140 1.020 3.685 1.250 ;
        RECT  2.910 1.020 3.140 2.835 ;
        RECT  2.745 2.605 2.910 2.835 ;
        RECT  2.515 2.605 2.745 3.455 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.620 6.315 1.965 ;
        RECT  5.740 1.620 6.020 2.375 ;
        RECT  4.340 2.135 5.740 2.375 ;
        RECT  3.370 1.770 4.340 2.375 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.470 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.260 -0.235 8.400 0.235 ;
        RECT  7.880 -0.235 8.260 0.465 ;
        RECT  5.285 -0.235 7.880 0.235 ;
        RECT  4.505 -0.235 5.285 0.465 ;
        RECT  2.085 -0.235 4.505 0.235 ;
        RECT  1.705 -0.235 2.085 1.180 ;
        RECT  0.625 -0.235 1.705 0.235 ;
        RECT  0.245 -0.235 0.625 0.940 ;
        RECT  0.000 -0.235 0.245 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.200 3.685 8.400 4.155 ;
        RECT  7.820 2.305 8.200 4.155 ;
        RECT  6.675 3.685 7.820 4.155 ;
        RECT  6.295 3.085 6.675 4.155 ;
        RECT  5.115 3.685 6.295 4.155 ;
        RECT  4.735 3.085 5.115 4.155 ;
        RECT  3.560 3.685 4.735 4.155 ;
        RECT  3.180 3.085 3.560 4.155 ;
        RECT  2.090 3.685 3.180 4.155 ;
        RECT  1.710 2.305 2.090 4.155 ;
        RECT  0.630 3.685 1.710 4.155 ;
        RECT  0.250 2.480 0.630 4.155 ;
        RECT  0.000 3.685 0.250 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.310 1.020 6.350 1.250 ;
        RECT  5.840 2.605 6.350 2.835 ;
        RECT  5.600 2.605 5.840 3.415 ;
        RECT  4.225 2.605 5.600 2.835 ;
        RECT  3.995 2.605 4.225 3.405 ;
        RECT  3.140 2.605 3.995 2.835 ;
        RECT  3.140 1.020 3.685 1.250 ;
        RECT  2.910 1.020 3.140 2.835 ;
        RECT  2.745 2.605 2.910 2.835 ;
        RECT  2.515 2.605 2.745 3.455 ;
        RECT  7.785 0.820 8.025 2.015 ;
        RECT  7.560 0.820 7.785 1.050 ;
        RECT  7.330 0.560 7.560 1.050 ;
        RECT  5.990 0.560 7.330 0.790 ;
        RECT  5.760 0.560 5.990 1.035 ;
        RECT  4.800 0.805 5.760 1.035 ;
        RECT  4.800 1.540 5.280 1.880 ;
        RECT  4.570 0.805 4.800 1.880 ;
        RECT  4.215 0.805 4.570 1.035 ;
        RECT  3.985 0.560 4.215 1.035 ;
        RECT  2.655 0.560 3.985 0.790 ;
        RECT  2.380 0.560 2.655 1.895 ;
        RECT  1.285 1.665 2.380 1.895 ;
        RECT  1.055 0.495 1.285 3.105 ;
    END
END IND2D4BWP7T

MACRO IND3D0BWP7T
    CLASS CORE ;
    FOREIGN IND3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9387 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.595 3.220 2.745 ;
        RECT  2.820 0.595 2.940 0.825 ;
        RECT  1.505 2.515 2.940 2.745 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.700 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.650 2.100 1.590 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.730 0.465 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 -0.235 3.360 0.235 ;
        RECT  0.880 -0.235 1.260 0.790 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 3.685 3.360 4.155 ;
        RECT  2.015 3.450 2.380 4.155 ;
        RECT  1.300 3.685 2.015 4.155 ;
        RECT  0.950 3.450 1.300 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.945 1.655 1.475 1.885 ;
        RECT  0.705 1.115 0.945 3.215 ;
        RECT  0.465 1.115 0.705 1.355 ;
        RECT  0.180 2.985 0.705 3.215 ;
        RECT  0.235 0.500 0.465 1.355 ;
    END
END IND3D0BWP7T

MACRO IND3D1BWP7T
    CLASS CORE ;
    FOREIGN IND3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.7597 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 0.660 3.170 0.890 ;
        RECT  2.895 2.380 3.135 3.330 ;
        RECT  2.660 2.380 2.895 2.745 ;
        RECT  2.420 0.660 2.660 2.745 ;
        RECT  1.505 2.380 2.420 2.745 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.210 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.3303 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.175 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.575 1.600 0.700 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 -0.235 3.360 0.235 ;
        RECT  0.920 -0.235 1.300 0.465 ;
        RECT  0.000 -0.235 0.920 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.420 3.685 3.360 4.155 ;
        RECT  2.055 3.450 2.420 4.155 ;
        RECT  1.090 3.685 2.055 4.155 ;
        RECT  0.740 3.450 1.090 4.155 ;
        RECT  0.000 3.685 0.740 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.265 0.705 1.495 1.970 ;
        RECT  0.530 0.705 1.265 0.940 ;
        RECT  0.345 2.510 0.540 2.750 ;
        RECT  0.345 0.470 0.530 0.940 ;
        RECT  0.115 0.470 0.345 2.750 ;
    END
END IND3D1BWP7T

MACRO IND3D2BWP7T
    CLASS CORE ;
    FOREIGN IND3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.8211 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.900 1.020 5.765 1.250 ;
        RECT  5.480 2.480 5.710 3.405 ;
        RECT  4.900 2.480 5.480 2.730 ;
        RECT  4.620 1.020 4.900 2.730 ;
        RECT  4.230 2.480 4.620 2.730 ;
        RECT  4.000 2.480 4.230 3.405 ;
        RECT  2.065 2.480 4.000 2.730 ;
        RECT  1.835 2.480 2.065 3.400 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.675 6.020 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.675 4.360 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.880 -0.235 6.720 0.235 ;
        RECT  2.500 -0.235 2.880 0.785 ;
        RECT  1.290 -0.235 2.500 0.235 ;
        RECT  0.930 -0.235 1.290 0.465 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.510 3.685 6.720 4.155 ;
        RECT  6.130 2.560 6.510 4.155 ;
        RECT  5.050 3.685 6.130 4.155 ;
        RECT  4.670 3.005 5.050 4.155 ;
        RECT  3.585 3.685 4.670 4.155 ;
        RECT  3.205 3.060 3.585 4.155 ;
        RECT  2.885 3.685 3.205 4.155 ;
        RECT  2.505 3.060 2.885 4.155 ;
        RECT  1.325 3.685 2.505 4.155 ;
        RECT  0.945 3.055 1.325 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.145 0.540 6.485 1.240 ;
        RECT  3.225 0.540 6.145 0.770 ;
        RECT  2.070 1.020 4.285 1.250 ;
        RECT  1.265 1.715 2.330 1.945 ;
        RECT  1.840 0.635 2.070 1.250 ;
        RECT  1.025 0.730 1.265 2.760 ;
        RECT  0.180 0.730 1.025 0.960 ;
        RECT  0.465 2.520 1.025 2.760 ;
        RECT  0.235 2.520 0.465 3.330 ;
    END
END IND3D2BWP7T

MACRO IND4D0BWP7T
    CLASS CORE ;
    FOREIGN IND4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9848 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 0.490 3.750 0.720 ;
        RECT  2.940 0.490 3.220 2.725 ;
        RECT  1.500 2.495 2.940 2.725 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 1.210 3.780 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.695 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.650 2.100 1.590 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.730 0.465 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 -0.235 3.920 0.235 ;
        RECT  0.880 -0.235 1.260 0.795 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 3.685 3.920 4.155 ;
        RECT  3.450 3.370 3.695 4.155 ;
        RECT  3.075 3.685 3.450 4.155 ;
        RECT  2.830 3.370 3.075 4.155 ;
        RECT  2.455 3.685 2.830 4.155 ;
        RECT  2.210 3.370 2.455 4.155 ;
        RECT  1.870 3.685 2.210 4.155 ;
        RECT  1.625 3.370 1.870 4.155 ;
        RECT  1.300 3.685 1.625 4.155 ;
        RECT  0.945 3.450 1.300 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.940 1.695 1.470 1.925 ;
        RECT  0.700 1.150 0.940 3.170 ;
        RECT  0.465 1.150 0.700 1.390 ;
        RECT  0.180 2.940 0.700 3.170 ;
        RECT  0.235 0.465 0.465 1.390 ;
    END
END IND4D0BWP7T

MACRO IND4D1BWP7T
    CLASS CORE ;
    FOREIGN IND4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.9896 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.945 0.495 4.175 1.345 ;
        RECT  3.780 1.105 3.945 1.345 ;
        RECT  3.500 1.105 3.780 2.795 ;
        RECT  3.425 2.565 3.500 2.795 ;
        RECT  3.195 2.565 3.425 3.375 ;
        RECT  1.985 2.565 3.195 2.795 ;
        RECT  1.755 2.565 1.985 3.375 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.610 4.340 2.710 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.650 3.220 1.830 ;
        RECT  2.655 1.600 2.940 1.830 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.170 2.180 2.190 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.295 -0.235 4.480 0.235 ;
        RECT  0.935 -0.235 1.295 0.470 ;
        RECT  0.000 -0.235 0.935 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.220 3.685 4.480 4.155 ;
        RECT  3.840 3.045 4.220 4.155 ;
        RECT  2.780 3.685 3.840 4.155 ;
        RECT  2.400 3.045 2.780 4.155 ;
        RECT  1.335 3.685 2.400 4.155 ;
        RECT  0.955 2.995 1.335 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.215 1.660 1.490 1.895 ;
        RECT  0.965 0.700 1.215 2.670 ;
        RECT  0.465 0.700 0.965 0.940 ;
        RECT  0.180 2.440 0.965 2.670 ;
        RECT  0.235 0.540 0.465 0.940 ;
    END
END IND4D1BWP7T

MACRO IND4D2BWP7T
    CLASS CORE ;
    FOREIGN IND4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.4664 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.160 1.005 7.500 1.440 ;
        RECT  7.215 2.580 7.445 3.415 ;
        RECT  7.140 2.580 7.215 2.820 ;
        RECT  7.140 1.210 7.160 1.440 ;
        RECT  6.860 1.210 7.140 2.820 ;
        RECT  6.005 2.580 6.860 2.820 ;
        RECT  5.775 2.580 6.005 3.410 ;
        RECT  3.865 2.580 5.775 2.820 ;
        RECT  3.635 2.580 3.865 3.410 ;
        RECT  2.425 2.580 3.635 2.820 ;
        RECT  2.195 2.580 2.425 3.410 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.740 1.770 8.260 2.150 ;
        RECT  7.400 1.680 7.740 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.8388 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.210 6.580 2.150 ;
        RECT  6.015 1.625 6.300 1.965 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8388 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 3.785 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 -0.235 8.400 0.235 ;
        RECT  2.175 -0.235 2.555 0.670 ;
        RECT  1.280 -0.235 2.175 0.235 ;
        RECT  0.940 -0.235 1.280 0.515 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.220 3.685 8.400 4.155 ;
        RECT  7.880 2.585 8.220 4.155 ;
        RECT  6.780 3.685 7.880 4.155 ;
        RECT  6.440 3.120 6.780 4.155 ;
        RECT  5.340 3.685 6.440 4.155 ;
        RECT  5.000 3.090 5.340 4.155 ;
        RECT  4.640 3.685 5.000 4.155 ;
        RECT  4.300 3.090 4.640 4.155 ;
        RECT  3.200 3.685 4.300 4.155 ;
        RECT  2.860 3.095 3.200 4.155 ;
        RECT  1.705 3.685 2.860 4.155 ;
        RECT  1.475 3.065 1.705 4.155 ;
        RECT  1.185 3.685 1.475 4.155 ;
        RECT  0.955 3.065 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.935 0.495 8.165 1.305 ;
        RECT  5.245 0.495 7.935 0.725 ;
        RECT  5.760 1.020 6.060 1.250 ;
        RECT  5.530 1.020 5.760 1.935 ;
        RECT  4.490 1.705 5.530 1.935 ;
        RECT  5.015 0.495 5.245 1.385 ;
        RECT  3.205 0.465 4.700 0.695 ;
        RECT  4.260 1.020 4.490 1.935 ;
        RECT  3.640 1.020 4.260 1.250 ;
        RECT  2.975 0.465 3.205 1.275 ;
        RECT  1.480 1.020 2.975 1.275 ;
        RECT  1.845 1.695 2.710 1.925 ;
        RECT  1.615 1.695 1.845 2.770 ;
        RECT  0.470 2.540 1.615 2.770 ;
        RECT  0.465 2.540 0.470 3.350 ;
        RECT  0.235 0.495 0.465 3.350 ;
    END
END IND4D2BWP7T

MACRO INR2D0BWP7T
    CLASS CORE ;
    FOREIGN INR2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.5988 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 3.040 2.620 3.270 ;
        RECT  1.820 0.915 2.100 3.270 ;
        RECT  1.560 0.915 1.820 1.145 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.770 2.660 2.710 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 -0.235 2.800 0.235 ;
        RECT  2.335 -0.235 2.575 1.200 ;
        RECT  0.000 -0.235 2.335 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 3.685 2.800 4.155 ;
        RECT  0.900 3.130 1.280 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.000 1.655 1.520 1.885 ;
        RECT  0.760 0.595 1.000 2.680 ;
        RECT  0.180 0.595 0.760 0.825 ;
        RECT  0.465 2.450 0.760 2.680 ;
        RECT  0.235 2.450 0.465 3.415 ;
    END
END INR2D0BWP7T

MACRO INR2D1BWP7T
    CLASS CORE ;
    FOREIGN INR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1976 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 3.030 2.640 3.270 ;
        RECT  1.850 1.170 2.100 3.270 ;
        RECT  1.820 0.495 1.850 3.270 ;
        RECT  1.610 0.495 1.820 1.450 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.645 2.660 2.710 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.470 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 -0.235 2.800 0.235 ;
        RECT  2.330 -0.235 2.575 1.310 ;
        RECT  0.520 -0.235 2.330 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 3.685 2.800 4.155 ;
        RECT  0.935 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.935 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.075 1.710 1.545 1.940 ;
        RECT  0.845 0.995 1.075 3.225 ;
        RECT  0.180 0.995 0.845 1.225 ;
        RECT  0.170 2.995 0.845 3.225 ;
    END
END INR2D1BWP7T

MACRO INR2D2BWP7T
    CLASS CORE ;
    FOREIGN INR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8746 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.295 0.690 3.525 1.310 ;
        RECT  3.220 1.050 3.295 1.310 ;
        RECT  2.940 1.050 3.220 2.815 ;
        RECT  2.045 1.050 2.940 1.310 ;
        RECT  2.500 2.585 2.940 2.815 ;
        RECT  1.815 0.690 2.045 1.310 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.660 2.660 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.730 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 1.195 ;
        RECT  2.875 -0.235 3.940 0.235 ;
        RECT  2.495 -0.235 2.875 0.785 ;
        RECT  1.355 -0.235 2.495 0.235 ;
        RECT  0.975 -0.235 1.355 0.800 ;
        RECT  0.000 -0.235 0.975 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 3.685 4.480 4.155 ;
        RECT  4.015 2.250 4.245 4.155 ;
        RECT  1.310 3.685 4.015 4.155 ;
        RECT  0.970 3.065 1.310 4.155 ;
        RECT  0.000 3.685 0.970 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.535 1.610 3.765 3.355 ;
        RECT  2.130 3.115 3.535 3.355 ;
        RECT  1.890 2.535 2.130 3.355 ;
        RECT  1.490 2.535 1.890 2.765 ;
        RECT  1.250 1.110 1.490 2.765 ;
        RECT  0.465 1.110 1.250 1.350 ;
        RECT  0.470 2.535 1.250 2.765 ;
        RECT  0.230 2.535 0.470 3.400 ;
        RECT  0.235 0.690 0.465 1.350 ;
    END
END INR2D2BWP7T

MACRO INR2D4BWP7T
    CLASS CORE ;
    FOREIGN INR2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.9273 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.550 0.725 7.450 2.765 ;
        RECT  2.450 0.725 6.550 0.955 ;
        RECT  3.215 2.535 6.550 2.765 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.620 6.315 1.965 ;
        RECT  5.740 1.620 6.020 2.305 ;
        RECT  3.780 2.065 5.740 2.305 ;
        RECT  2.940 1.770 3.780 2.305 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.470 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.220 -0.235 8.400 0.235 ;
        RECT  7.880 -0.235 8.220 1.140 ;
        RECT  6.650 -0.235 7.880 0.235 ;
        RECT  6.310 -0.235 6.650 0.465 ;
        RECT  5.090 -0.235 6.310 0.235 ;
        RECT  4.750 -0.235 5.090 0.465 ;
        RECT  3.550 -0.235 4.750 0.235 ;
        RECT  3.210 -0.235 3.550 0.465 ;
        RECT  2.085 -0.235 3.210 0.235 ;
        RECT  1.705 -0.235 2.085 1.180 ;
        RECT  0.625 -0.235 1.705 0.235 ;
        RECT  0.245 -0.235 0.625 0.940 ;
        RECT  0.000 -0.235 0.245 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.220 3.685 8.400 4.155 ;
        RECT  7.880 3.455 8.220 4.155 ;
        RECT  5.115 3.685 7.880 4.155 ;
        RECT  4.735 3.455 5.115 4.155 ;
        RECT  2.090 3.685 4.735 4.155 ;
        RECT  1.710 2.480 2.090 4.155 ;
        RECT  0.630 3.685 1.710 4.155 ;
        RECT  0.250 2.480 0.630 4.155 ;
        RECT  0.000 3.685 0.250 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.450 0.725 6.350 0.955 ;
        RECT  3.215 2.535 6.350 2.765 ;
        RECT  7.680 1.620 7.910 3.225 ;
        RECT  2.655 2.995 7.680 3.225 ;
        RECT  4.745 1.585 5.320 1.815 ;
        RECT  4.510 1.250 4.745 1.815 ;
        RECT  2.655 1.250 4.510 1.480 ;
        RECT  2.425 1.250 2.655 3.225 ;
        RECT  1.285 1.665 2.425 1.895 ;
        RECT  1.055 0.465 1.285 3.375 ;
    END
END INR2D4BWP7T

MACRO INR2XD0BWP7T
    CLASS CORE ;
    FOREIGN INR2XD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9276 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 3.040 2.620 3.270 ;
        RECT  1.820 0.915 2.100 3.270 ;
        RECT  1.560 0.915 1.820 1.145 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.615 2.660 2.710 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 -0.235 2.800 0.235 ;
        RECT  2.335 -0.235 2.610 1.200 ;
        RECT  0.000 -0.235 2.335 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 3.685 2.800 4.155 ;
        RECT  0.900 3.105 1.280 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.000 1.655 1.520 1.885 ;
        RECT  0.760 0.635 1.000 2.680 ;
        RECT  0.180 0.635 0.760 0.865 ;
        RECT  0.465 2.450 0.760 2.680 ;
        RECT  0.235 2.450 0.465 3.390 ;
    END
END INR2XD0BWP7T

MACRO INR2XD1BWP7T
    CLASS CORE ;
    FOREIGN INR2XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.4548 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 2.525 2.860 2.755 ;
        RECT  2.150 0.965 2.380 1.645 ;
        RECT  2.120 1.415 2.150 1.645 ;
        RECT  1.820 1.415 2.120 2.755 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 1.770 3.780 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 -0.235 4.480 0.235 ;
        RECT  3.070 -0.235 3.300 0.780 ;
        RECT  1.460 -0.235 3.070 0.235 ;
        RECT  1.230 -0.235 1.460 0.725 ;
        RECT  0.000 -0.235 1.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 3.685 4.480 4.155 ;
        RECT  3.940 2.570 4.320 4.155 ;
        RECT  1.440 3.685 3.940 4.155 ;
        RECT  1.060 2.970 1.440 4.155 ;
        RECT  0.000 3.685 1.060 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.010 1.125 4.240 1.975 ;
        RECT  2.840 1.125 4.010 1.355 ;
        RECT  3.240 2.475 3.580 3.220 ;
        RECT  1.800 2.990 3.240 3.220 ;
        RECT  2.610 0.465 2.840 1.355 ;
        RECT  1.920 0.465 2.610 0.695 ;
        RECT  1.690 0.465 1.920 1.185 ;
        RECT  0.960 0.955 1.690 1.185 ;
        RECT  0.960 1.670 1.520 1.900 ;
        RECT  0.910 0.650 0.960 1.900 ;
        RECT  0.680 0.650 0.910 2.710 ;
        RECT  0.200 0.650 0.680 0.890 ;
        RECT  0.485 2.470 0.680 2.710 ;
        RECT  0.255 2.470 0.485 3.365 ;
    END
END INR2XD1BWP7T

MACRO INR2XD2BWP7T
    CLASS CORE ;
    FOREIGN INR2XD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0946 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.770 0.965 5.005 2.660 ;
        RECT  2.245 2.380 4.770 2.660 ;
        RECT  2.015 0.965 2.245 2.660 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.305 1.600 4.535 2.100 ;
        RECT  2.715 1.770 4.305 2.100 ;
        RECT  2.485 1.595 2.715 2.100 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.670 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 -0.235 6.160 0.235 ;
        RECT  5.695 -0.235 5.925 0.725 ;
        RECT  4.080 -0.235 5.695 0.235 ;
        RECT  3.850 -0.235 4.080 0.820 ;
        RECT  3.165 -0.235 3.850 0.235 ;
        RECT  2.935 -0.235 3.165 0.820 ;
        RECT  1.315 -0.235 2.935 0.235 ;
        RECT  1.085 -0.235 1.315 0.810 ;
        RECT  0.000 -0.235 1.085 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.000 3.685 6.160 4.155 ;
        RECT  5.620 2.305 6.000 4.155 ;
        RECT  3.700 3.685 5.620 4.155 ;
        RECT  3.320 2.950 3.700 4.155 ;
        RECT  1.260 3.685 3.320 4.155 ;
        RECT  0.880 2.950 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.465 1.600 5.695 1.980 ;
        RECT  5.235 0.465 5.465 1.980 ;
        RECT  4.540 0.465 5.235 0.695 ;
        RECT  4.310 0.465 4.540 1.280 ;
        RECT  3.850 1.050 4.310 1.280 ;
        RECT  3.200 1.050 3.850 1.540 ;
        RECT  2.705 1.050 3.200 1.280 ;
        RECT  2.475 0.465 2.705 1.280 ;
        RECT  1.775 0.465 2.475 0.695 ;
        RECT  1.560 0.465 1.775 1.300 ;
        RECT  1.545 0.465 1.560 2.710 ;
        RECT  1.320 1.070 1.545 2.710 ;
        RECT  0.465 1.070 1.320 1.300 ;
        RECT  0.465 2.470 1.320 2.710 ;
        RECT  0.235 0.465 0.465 1.300 ;
        RECT  0.235 2.470 0.465 3.390 ;
    END
END INR2XD2BWP7T

MACRO INR2XD4BWP7T
    CLASS CORE ;
    FOREIGN INR2XD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.2330 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.890 2.335 10.545 2.710 ;
        RECT  9.595 0.520 9.825 1.320 ;
        RECT  8.385 0.970 9.595 1.320 ;
        RECT  8.155 0.525 8.385 1.320 ;
        RECT  6.945 0.970 8.155 1.320 ;
        RECT  6.890 0.525 6.945 1.320 ;
        RECT  6.715 0.525 6.890 2.710 ;
        RECT  5.990 0.970 6.715 2.710 ;
        RECT  5.505 0.970 5.990 1.320 ;
        RECT  5.275 0.525 5.505 1.320 ;
        RECT  4.065 0.970 5.275 1.320 ;
        RECT  3.835 0.525 4.065 1.320 ;
        RECT  2.625 0.970 3.835 1.320 ;
        RECT  2.395 0.525 2.625 1.320 ;
        RECT  1.185 0.970 2.395 1.320 ;
        RECT  0.955 0.525 1.185 1.320 ;
        END
    END ZN
    PIN B1
        ANTENNAGATEAREA 2.6442 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 1.595 4.925 1.825 ;
        RECT  2.360 1.595 3.240 2.150 ;
        RECT  0.660 1.595 2.360 1.825 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.415 1.210 12.740 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.720 -0.235 12.880 0.235 ;
        RECT  12.340 -0.235 12.720 0.890 ;
        RECT  11.210 -0.235 12.340 0.235 ;
        RECT  10.970 -0.235 11.210 1.335 ;
        RECT  10.660 -0.235 10.970 0.235 ;
        RECT  10.390 -0.235 10.660 0.815 ;
        RECT  9.160 -0.235 10.390 0.235 ;
        RECT  8.820 -0.235 9.160 0.670 ;
        RECT  7.720 -0.235 8.820 0.235 ;
        RECT  7.380 -0.235 7.720 0.670 ;
        RECT  6.280 -0.235 7.380 0.235 ;
        RECT  5.940 -0.235 6.280 0.670 ;
        RECT  4.840 -0.235 5.940 0.235 ;
        RECT  4.500 -0.235 4.840 0.670 ;
        RECT  3.400 -0.235 4.500 0.235 ;
        RECT  3.060 -0.235 3.400 0.670 ;
        RECT  1.960 -0.235 3.060 0.235 ;
        RECT  1.620 -0.235 1.960 0.670 ;
        RECT  0.520 -0.235 1.620 0.235 ;
        RECT  0.180 -0.235 0.520 0.745 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.720 3.685 12.880 4.155 ;
        RECT  12.340 2.565 12.720 4.155 ;
        RECT  11.275 3.685 12.340 4.155 ;
        RECT  10.895 3.190 11.275 4.155 ;
        RECT  4.860 3.685 10.895 4.155 ;
        RECT  4.480 3.090 4.860 4.155 ;
        RECT  3.420 3.685 4.480 4.155 ;
        RECT  3.040 3.090 3.420 4.155 ;
        RECT  1.980 3.685 3.040 4.155 ;
        RECT  1.600 3.090 1.980 4.155 ;
        RECT  0.540 3.685 1.600 4.155 ;
        RECT  0.160 2.570 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.090 2.335 10.545 2.710 ;
        RECT  9.595 0.520 9.825 1.320 ;
        RECT  8.385 0.970 9.595 1.320 ;
        RECT  8.155 0.525 8.385 1.320 ;
        RECT  7.090 0.970 8.155 1.320 ;
        RECT  5.505 0.970 5.790 1.320 ;
        RECT  5.275 0.525 5.505 1.320 ;
        RECT  4.065 0.970 5.275 1.320 ;
        RECT  3.835 0.525 4.065 1.320 ;
        RECT  2.625 0.970 3.835 1.320 ;
        RECT  2.395 0.525 2.625 1.320 ;
        RECT  1.185 0.970 2.395 1.320 ;
        RECT  0.955 0.525 1.185 1.320 ;
        RECT  11.695 0.495 11.925 3.430 ;
        RECT  7.460 1.595 11.695 1.825 ;
        RECT  5.505 2.950 9.880 3.180 ;
        RECT  5.275 2.170 5.505 3.450 ;
        RECT  4.065 2.470 5.275 2.760 ;
        RECT  3.835 2.470 4.065 3.410 ;
        RECT  2.625 2.470 3.835 2.760 ;
        RECT  2.395 2.470 2.625 3.410 ;
        RECT  1.185 2.470 2.395 2.760 ;
        RECT  0.955 2.470 1.185 3.410 ;
    END
END INR2XD4BWP7T

MACRO INR3D0BWP7T
    CLASS CORE ;
    FOREIGN INR3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2176 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 0.580 3.780 3.360 ;
        RECT  1.960 3.130 3.455 3.360 ;
        RECT  1.725 0.560 1.960 3.360 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.665 2.660 2.750 ;
        RECT  2.200 1.665 2.380 1.895 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.920 -0.235 3.920 0.235 ;
        RECT  2.540 -0.235 2.920 0.855 ;
        RECT  1.260 -0.235 2.540 0.235 ;
        RECT  0.880 -0.235 1.260 0.825 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.360 3.685 3.920 4.155 ;
        RECT  0.980 3.050 1.360 4.155 ;
        RECT  0.000 3.685 0.980 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.255 1.600 1.485 2.795 ;
        RECT  0.355 2.565 1.255 2.795 ;
        RECT  0.355 0.595 0.520 0.825 ;
        RECT  0.115 0.595 0.355 2.795 ;
    END
END INR3D0BWP7T

MACRO INR3D1BWP7T
    CLASS CORE ;
    FOREIGN INR3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.6724 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 0.700 4.315 2.245 ;
        RECT  1.670 0.700 4.085 0.980 ;
        RECT  3.780 2.015 4.085 2.245 ;
        RECT  3.500 2.015 3.780 2.790 ;
        RECT  2.705 2.560 3.500 2.790 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.6282 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.6282 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.625 1.210 3.855 1.745 ;
        RECT  2.145 1.210 3.625 1.450 ;
        RECT  1.820 1.210 2.145 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.575 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 -0.235 5.040 0.235 ;
        RECT  2.430 -0.235 2.770 0.465 ;
        RECT  1.290 -0.235 2.430 0.235 ;
        RECT  0.910 -0.235 1.290 0.765 ;
        RECT  0.000 -0.235 0.910 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 3.685 5.040 4.155 ;
        RECT  4.575 3.010 4.805 4.155 ;
        RECT  1.185 3.685 4.575 4.155 ;
        RECT  0.955 3.195 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.545 1.565 4.775 2.780 ;
        RECT  4.345 2.550 4.545 2.780 ;
        RECT  4.115 2.550 4.345 3.250 ;
        RECT  2.265 3.020 4.115 3.250 ;
        RECT  2.035 2.545 2.265 3.250 ;
        RECT  1.475 2.545 2.035 2.775 ;
        RECT  1.245 1.660 1.475 2.775 ;
        RECT  0.465 2.540 1.245 2.775 ;
        RECT  0.345 0.595 0.540 0.980 ;
        RECT  0.345 2.540 0.465 3.440 ;
        RECT  0.115 0.595 0.345 3.440 ;
    END
END INR3D1BWP7T

MACRO INR3D2BWP7T
    CLASS CORE ;
    FOREIGN INR3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.4072 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.485 0.465 5.720 1.310 ;
        RECT  5.485 2.000 5.715 2.910 ;
        RECT  4.900 1.020 5.485 1.310 ;
        RECT  4.900 2.000 5.485 2.280 ;
        RECT  4.620 1.020 4.900 2.280 ;
        RECT  4.245 1.020 4.620 1.310 ;
        RECT  4.015 0.465 4.245 1.310 ;
        RECT  2.065 1.020 4.015 1.310 ;
        RECT  1.835 0.465 2.065 1.310 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.255 1.660 6.580 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 4.340 2.150 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 -0.235 6.720 0.235 ;
        RECT  6.180 -0.235 6.560 1.200 ;
        RECT  5.040 -0.235 6.180 0.235 ;
        RECT  4.660 -0.235 5.040 0.790 ;
        RECT  3.600 -0.235 4.660 0.235 ;
        RECT  3.220 -0.235 3.600 0.790 ;
        RECT  2.900 -0.235 3.220 0.235 ;
        RECT  2.520 -0.235 2.900 0.790 ;
        RECT  1.350 -0.235 2.520 0.235 ;
        RECT  0.970 -0.235 1.350 0.965 ;
        RECT  0.000 -0.235 0.970 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.880 3.685 6.720 4.155 ;
        RECT  2.540 3.455 2.880 4.155 ;
        RECT  1.340 3.685 2.540 4.155 ;
        RECT  0.960 3.000 1.340 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.255 3.040 6.485 3.455 ;
        RECT  4.965 3.215 6.255 3.455 ;
        RECT  4.735 2.510 4.965 3.455 ;
        RECT  3.240 2.510 4.735 2.740 ;
        RECT  2.065 2.985 4.300 3.225 ;
        RECT  1.530 1.685 2.360 1.915 ;
        RECT  1.835 2.415 2.065 3.225 ;
        RECT  1.300 1.685 1.530 2.720 ;
        RECT  0.465 2.490 1.300 2.720 ;
        RECT  0.235 0.465 0.465 3.350 ;
    END
END INR3D2BWP7T

MACRO INR4D0BWP7T
    CLASS CORE ;
    FOREIGN INR4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.3572 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.000 4.340 3.360 ;
        RECT  3.710 1.000 4.060 1.230 ;
        RECT  3.975 2.935 4.060 3.360 ;
        RECT  1.960 3.130 3.975 3.360 ;
        RECT  3.480 0.480 3.710 1.230 ;
        RECT  3.230 0.480 3.480 0.710 ;
        RECT  1.725 0.465 1.960 3.360 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.670 3.830 2.710 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.025 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.665 2.660 2.750 ;
        RECT  2.200 1.665 2.380 1.895 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.585 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 -0.235 4.480 0.235 ;
        RECT  3.940 -0.235 4.320 0.720 ;
        RECT  2.840 -0.235 3.940 0.235 ;
        RECT  2.460 -0.235 2.840 0.710 ;
        RECT  1.195 -0.235 2.460 0.235 ;
        RECT  0.945 -0.235 1.195 0.810 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.360 3.685 4.480 4.155 ;
        RECT  0.980 3.050 1.360 4.155 ;
        RECT  0.000 3.685 0.980 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.255 1.600 1.485 2.795 ;
        RECT  0.355 2.565 1.255 2.795 ;
        RECT  0.355 0.520 0.520 0.750 ;
        RECT  0.115 0.520 0.355 2.795 ;
    END
END INR4D0BWP7T

MACRO INR4D1BWP7T
    CLASS CORE ;
    FOREIGN INR4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.4958 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 2.380 4.050 2.660 ;
        RECT  3.565 0.595 3.795 0.935 ;
        RECT  2.885 0.695 3.565 0.935 ;
        RECT  2.655 0.695 2.885 2.660 ;
        RECT  1.185 0.695 2.655 0.925 ;
        RECT  0.955 0.585 1.185 0.925 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.6192 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 4.340 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.6192 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.425 1.210 1.590 1.590 ;
        RECT  1.195 1.210 1.425 1.825 ;
        RECT  0.700 1.210 1.195 1.590 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.6192 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.220 2.375 2.340 ;
        RECT  0.465 2.100 2.145 2.340 ;
        RECT  0.140 1.210 0.465 2.340 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.295 -0.235 6.720 0.235 ;
        RECT  5.955 -0.235 6.295 0.785 ;
        RECT  4.570 -0.235 5.955 0.235 ;
        RECT  4.230 -0.235 4.570 0.880 ;
        RECT  3.090 -0.235 4.230 0.235 ;
        RECT  2.750 -0.235 3.090 0.465 ;
        RECT  2.000 -0.235 2.750 0.235 ;
        RECT  1.660 -0.235 2.000 0.465 ;
        RECT  0.520 -0.235 1.660 0.235 ;
        RECT  0.180 -0.235 0.520 0.670 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.540 3.685 6.720 4.155 ;
        RECT  6.200 2.490 6.540 4.155 ;
        RECT  1.750 3.685 6.200 4.155 ;
        RECT  1.370 3.140 1.750 4.155 ;
        RECT  0.000 3.685 1.370 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.185 2.395 5.820 2.625 ;
        RECT  5.185 0.575 5.575 0.805 ;
        RECT  2.280 3.225 5.205 3.455 ;
        RECT  4.955 0.575 5.185 2.625 ;
        RECT  3.130 1.240 4.955 1.470 ;
        RECT  2.050 2.645 2.280 3.455 ;
        RECT  0.465 2.645 2.050 2.875 ;
        RECT  0.235 2.645 0.465 3.455 ;
    END
END INR4D1BWP7T

MACRO INR4D2BWP7T
    CLASS CORE ;
    FOREIGN INR4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.6396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.180 2.580 13.660 2.810 ;
        RECT  12.655 0.475 12.885 1.370 ;
        RECT  12.180 1.140 12.655 1.370 ;
        RECT  11.880 1.140 12.180 2.810 ;
        RECT  10.005 1.140 11.880 1.370 ;
        RECT  9.775 0.475 10.005 1.370 ;
        RECT  6.205 1.140 9.775 1.370 ;
        RECT  5.975 0.475 6.205 1.370 ;
        RECT  3.325 1.140 5.975 1.370 ;
        RECT  3.095 0.475 3.325 1.370 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.580 1.630 14.420 2.150 ;
        RECT  12.470 1.630 13.580 1.860 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.500 1.630 10.930 1.860 ;
        RECT  9.660 1.630 10.500 2.150 ;
        RECT  8.915 1.630 9.660 1.860 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.580 1.630 6.975 1.860 ;
        RECT  5.740 1.630 6.580 2.150 ;
        RECT  4.960 1.630 5.740 1.860 ;
        END
    END B1
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.700 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.700 1.195 ;
        RECT  12.220 -0.235 13.320 0.235 ;
        RECT  11.840 -0.235 12.220 0.890 ;
        RECT  10.830 -0.235 11.840 0.235 ;
        RECT  10.450 -0.235 10.830 0.890 ;
        RECT  9.340 -0.235 10.450 0.235 ;
        RECT  8.960 -0.235 9.340 0.890 ;
        RECT  7.030 -0.235 8.960 0.235 ;
        RECT  6.650 -0.235 7.030 0.890 ;
        RECT  5.540 -0.235 6.650 0.235 ;
        RECT  5.160 -0.235 5.540 0.890 ;
        RECT  4.150 -0.235 5.160 0.235 ;
        RECT  3.770 -0.235 4.150 0.890 ;
        RECT  2.660 -0.235 3.770 0.235 ;
        RECT  2.280 -0.235 2.660 1.195 ;
        RECT  0.540 -0.235 2.280 0.235 ;
        RECT  0.160 -0.235 0.540 0.850 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.120 3.685 14.560 4.155 ;
        RECT  3.740 2.630 4.120 4.155 ;
        RECT  2.680 3.685 3.740 4.155 ;
        RECT  2.300 2.630 2.680 4.155 ;
        RECT  0.540 3.685 2.300 4.155 ;
        RECT  0.160 2.535 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.040 2.635 14.380 3.385 ;
        RECT  11.445 3.155 14.040 3.385 ;
        RECT  11.215 2.380 11.445 3.385 ;
        RECT  10.005 2.380 11.215 2.610 ;
        RECT  10.495 2.900 10.725 3.455 ;
        RECT  9.285 3.225 10.495 3.455 ;
        RECT  9.775 2.380 10.005 2.965 ;
        RECT  8.565 2.380 9.775 2.610 ;
        RECT  9.055 2.900 9.285 3.455 ;
        RECT  6.925 3.225 9.055 3.455 ;
        RECT  8.335 2.380 8.565 2.965 ;
        RECT  7.415 2.380 7.645 2.965 ;
        RECT  6.205 2.380 7.415 2.610 ;
        RECT  6.695 2.900 6.925 3.455 ;
        RECT  5.485 3.225 6.695 3.455 ;
        RECT  5.975 2.380 6.205 2.965 ;
        RECT  4.765 2.380 5.975 2.610 ;
        RECT  5.255 2.900 5.485 3.455 ;
        RECT  4.535 2.105 4.765 3.385 ;
        RECT  3.325 2.105 4.535 2.345 ;
        RECT  1.185 1.630 4.240 1.860 ;
        RECT  3.095 2.105 3.325 3.385 ;
        RECT  1.885 2.105 3.095 2.345 ;
        RECT  1.650 2.105 1.885 3.380 ;
        RECT  0.955 0.475 1.185 3.380 ;
    END
END INR4D2BWP7T

MACRO INVD0BWP7T
    CLASS CORE ;
    FOREIGN INVD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6162 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 0.685 1.540 3.035 ;
        RECT  1.135 0.685 1.260 0.935 ;
        RECT  1.140 2.795 1.260 3.035 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.530 -0.235 1.680 0.235 ;
        RECT  0.290 -0.235 0.530 0.980 ;
        RECT  0.000 -0.235 0.290 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 3.685 1.680 4.155 ;
        RECT  0.300 2.750 0.540 4.155 ;
        RECT  0.000 3.685 0.300 4.155 ;
        END
    END VDD
END INVD0BWP7T

MACRO INVD10BWP7T
    CLASS CORE ;
    FOREIGN INVD10BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 6.3990 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.965 0.695 7.195 1.400 ;
        RECT  6.965 2.150 7.195 3.385 ;
        RECT  5.715 1.000 6.965 1.400 ;
        RECT  5.715 2.150 6.965 2.550 ;
        RECT  5.485 0.695 5.715 1.400 ;
        RECT  5.485 2.150 5.715 3.385 ;
        RECT  5.210 1.000 5.485 1.400 ;
        RECT  5.210 2.150 5.485 2.550 ;
        RECT  4.215 1.000 5.210 2.550 ;
        RECT  3.985 0.695 4.215 3.385 ;
        RECT  3.750 1.000 3.985 2.550 ;
        RECT  2.715 1.000 3.750 1.400 ;
        RECT  2.715 2.150 3.750 2.550 ;
        RECT  2.485 0.695 2.715 1.400 ;
        RECT  2.485 2.150 2.715 3.385 ;
        RECT  1.215 1.000 2.485 1.400 ;
        RECT  1.215 2.150 2.485 2.550 ;
        RECT  0.985 0.695 1.215 1.400 ;
        RECT  0.985 2.150 1.215 3.385 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 4.2660 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.630 3.215 1.920 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.010 -0.235 8.400 0.235 ;
        RECT  7.630 -0.235 8.010 1.195 ;
        RECT  6.530 -0.235 7.630 0.235 ;
        RECT  6.150 -0.235 6.530 0.765 ;
        RECT  5.050 -0.235 6.150 0.235 ;
        RECT  4.670 -0.235 5.050 0.765 ;
        RECT  3.550 -0.235 4.670 0.235 ;
        RECT  3.170 -0.235 3.550 0.770 ;
        RECT  2.055 -0.235 3.170 0.235 ;
        RECT  1.675 -0.235 2.055 0.770 ;
        RECT  0.540 -0.235 1.675 0.235 ;
        RECT  0.160 -0.235 0.540 0.945 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.010 3.685 8.400 4.155 ;
        RECT  7.630 2.305 8.010 4.155 ;
        RECT  6.530 3.685 7.630 4.155 ;
        RECT  6.150 2.780 6.530 4.155 ;
        RECT  5.050 3.685 6.150 4.155 ;
        RECT  4.670 2.780 5.050 4.155 ;
        RECT  3.550 3.685 4.670 4.155 ;
        RECT  3.170 2.780 3.550 4.155 ;
        RECT  2.055 3.685 3.170 4.155 ;
        RECT  1.675 2.780 2.055 4.155 ;
        RECT  0.570 3.685 1.675 4.155 ;
        RECT  0.190 2.595 0.570 4.155 ;
        RECT  0.000 3.685 0.190 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.965 0.695 7.195 1.400 ;
        RECT  6.965 2.150 7.195 3.385 ;
        RECT  5.715 1.000 6.965 1.400 ;
        RECT  5.715 2.150 6.965 2.550 ;
        RECT  5.485 0.695 5.715 1.400 ;
        RECT  5.485 2.150 5.715 3.385 ;
        RECT  5.410 1.000 5.485 1.400 ;
        RECT  5.410 2.150 5.485 2.550 ;
        RECT  2.715 1.000 3.550 1.400 ;
        RECT  2.715 2.150 3.550 2.550 ;
        RECT  2.485 0.695 2.715 1.400 ;
        RECT  2.485 2.150 2.715 3.385 ;
        RECT  1.215 1.000 2.485 1.400 ;
        RECT  1.215 2.150 2.485 2.550 ;
        RECT  0.985 0.695 1.215 1.400 ;
        RECT  0.985 2.150 1.215 3.385 ;
    END
END INVD10BWP7T

MACRO INVD12BWP7T
    CLASS CORE ;
    FOREIGN INVD12BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 7.7736 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.170 0.500 8.510 1.410 ;
        RECT  8.170 2.120 8.510 3.380 ;
        RECT  7.070 1.010 8.170 1.410 ;
        RECT  7.070 2.120 8.170 2.520 ;
        RECT  6.730 0.500 7.070 1.410 ;
        RECT  6.730 2.120 7.070 3.380 ;
        RECT  5.770 1.010 6.730 1.410 ;
        RECT  5.770 2.120 6.730 2.520 ;
        RECT  5.590 1.010 5.770 2.520 ;
        RECT  5.250 0.500 5.590 3.380 ;
        RECT  4.310 1.010 5.250 2.520 ;
        RECT  4.140 1.010 4.310 1.410 ;
        RECT  4.140 2.120 4.310 2.520 ;
        RECT  3.800 0.500 4.140 1.410 ;
        RECT  3.800 2.120 4.140 3.380 ;
        RECT  2.680 1.010 3.800 1.410 ;
        RECT  2.680 2.120 3.800 2.520 ;
        RECT  2.340 0.500 2.680 1.410 ;
        RECT  2.340 2.120 2.680 3.380 ;
        RECT  1.240 1.010 2.340 1.410 ;
        RECT  1.240 2.120 2.340 2.520 ;
        RECT  0.900 0.500 1.240 1.410 ;
        RECT  0.900 2.120 1.240 3.380 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 5.1192 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.640 3.940 1.890 ;
        RECT  0.135 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.270 -0.235 9.520 0.235 ;
        RECT  8.930 -0.235 9.270 1.195 ;
        RECT  7.790 -0.235 8.930 0.235 ;
        RECT  7.450 -0.235 7.790 0.760 ;
        RECT  6.310 -0.235 7.450 0.235 ;
        RECT  5.970 -0.235 6.310 0.760 ;
        RECT  4.860 -0.235 5.970 0.235 ;
        RECT  4.520 -0.235 4.860 0.760 ;
        RECT  3.400 -0.235 4.520 0.235 ;
        RECT  3.060 -0.235 3.400 0.760 ;
        RECT  1.960 -0.235 3.060 0.235 ;
        RECT  1.620 -0.235 1.960 0.760 ;
        RECT  0.520 -0.235 1.620 0.235 ;
        RECT  0.180 -0.235 0.520 0.910 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.270 3.685 9.520 4.155 ;
        RECT  8.930 2.305 9.270 4.155 ;
        RECT  7.790 3.685 8.930 4.155 ;
        RECT  7.450 2.750 7.790 4.155 ;
        RECT  6.310 3.685 7.450 4.155 ;
        RECT  5.970 2.750 6.310 4.155 ;
        RECT  4.860 3.685 5.970 4.155 ;
        RECT  4.520 2.750 4.860 4.155 ;
        RECT  3.400 3.685 4.520 4.155 ;
        RECT  3.060 2.750 3.400 4.155 ;
        RECT  1.960 3.685 3.060 4.155 ;
        RECT  1.620 2.750 1.960 4.155 ;
        RECT  0.520 3.685 1.620 4.155 ;
        RECT  0.180 2.510 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.170 0.500 8.510 1.410 ;
        RECT  8.170 2.120 8.510 3.380 ;
        RECT  7.070 1.010 8.170 1.410 ;
        RECT  7.070 2.120 8.170 2.520 ;
        RECT  6.730 0.500 7.070 1.410 ;
        RECT  6.730 2.120 7.070 3.380 ;
        RECT  5.970 1.010 6.730 1.410 ;
        RECT  5.970 2.120 6.730 2.520 ;
        RECT  3.800 0.500 4.110 1.410 ;
        RECT  3.800 2.120 4.110 3.380 ;
        RECT  2.680 1.010 3.800 1.410 ;
        RECT  2.680 2.120 3.800 2.520 ;
        RECT  2.340 0.500 2.680 1.410 ;
        RECT  2.340 2.120 2.680 3.380 ;
        RECT  1.240 1.010 2.340 1.410 ;
        RECT  1.240 2.120 2.340 2.520 ;
        RECT  0.900 0.500 1.240 1.410 ;
        RECT  0.900 2.120 1.240 3.380 ;
    END
END INVD12BWP7T

MACRO INVD1BWP7T
    CLASS CORE ;
    FOREIGN INVD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2324 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 0.475 1.540 3.380 ;
        RECT  1.160 0.475 1.260 1.205 ;
        RECT  1.160 2.290 1.260 3.380 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.605 0.925 1.945 ;
        RECT  0.135 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.580 -0.235 1.680 0.235 ;
        RECT  0.240 -0.235 0.580 0.890 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.590 3.685 1.680 4.155 ;
        RECT  0.250 2.515 0.590 4.155 ;
        RECT  0.000 3.685 0.250 4.155 ;
        END
    END VDD
END INVD1BWP7T

MACRO INVD1P5BWP7T
    CLASS CORE ;
    FOREIGN INVD1P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2679 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.070 1.540 2.710 ;
        RECT  1.235 1.070 1.260 1.300 ;
        RECT  1.235 2.330 1.260 2.710 ;
        RECT  1.005 0.630 1.235 1.300 ;
        RECT  1.005 2.330 1.235 3.415 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.6399 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.615 1.000 1.955 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.080 0.710 ;
        RECT  0.540 -0.235 1.700 0.235 ;
        RECT  0.160 -0.235 0.540 0.845 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 3.685 2.240 4.155 ;
        RECT  1.700 3.115 2.080 4.155 ;
        RECT  0.540 3.685 1.700 4.155 ;
        RECT  0.160 2.595 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
END INVD1P5BWP7T

MACRO INVD2BWP7T
    CLASS CORE ;
    FOREIGN INVD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 1.165 1.540 2.710 ;
        RECT  1.260 0.490 1.290 2.710 ;
        RECT  0.950 0.490 1.260 1.395 ;
        RECT  1.235 2.345 1.260 2.710 ;
        RECT  1.005 2.345 1.235 3.425 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.660 0.935 1.890 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 -0.235 2.240 0.235 ;
        RECT  1.775 -0.235 2.015 1.195 ;
        RECT  0.540 -0.235 1.775 0.235 ;
        RECT  0.160 -0.235 0.540 0.845 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.010 3.685 2.240 4.155 ;
        RECT  1.775 2.245 2.010 4.155 ;
        RECT  0.540 3.685 1.775 4.155 ;
        RECT  0.160 2.595 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
END INVD2BWP7T

MACRO INVD2P5BWP7T
    CLASS CORE ;
    FOREIGN INVD2P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.1490 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.075 2.660 2.655 ;
        RECT  1.910 1.075 2.380 1.310 ;
        RECT  0.470 2.425 2.380 2.655 ;
        RECT  1.665 0.895 1.910 1.310 ;
        RECT  0.475 1.075 1.665 1.310 ;
        RECT  0.230 0.465 0.475 1.310 ;
        RECT  0.230 2.425 0.470 3.355 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.0602 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.660 2.085 1.890 ;
        RECT  0.140 1.660 0.980 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 -0.235 2.800 0.235 ;
        RECT  2.325 -0.235 2.570 0.535 ;
        RECT  1.260 -0.235 2.325 0.235 ;
        RECT  0.900 -0.235 1.260 0.810 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 3.685 2.800 4.155 ;
        RECT  2.320 3.230 2.575 4.155 ;
        RECT  1.250 3.685 2.320 4.155 ;
        RECT  0.885 2.935 1.250 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
END INVD2P5BWP7T

MACRO INVD3BWP7T
    CLASS CORE ;
    FOREIGN INVD3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.4648 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.490 3.170 1.395 ;
        RECT  2.970 2.145 3.100 3.355 ;
        RECT  2.870 0.490 2.970 3.355 ;
        RECT  2.805 0.490 2.870 2.495 ;
        RECT  2.070 1.045 2.805 2.495 ;
        RECT  1.505 1.045 2.070 1.395 ;
        RECT  1.450 2.145 2.070 2.495 ;
        RECT  1.160 0.495 1.505 1.395 ;
        RECT  1.220 2.145 1.450 3.355 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.655 1.525 1.895 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 -0.235 3.360 0.235 ;
        RECT  1.970 -0.235 2.350 0.760 ;
        RECT  0.685 -0.235 1.970 0.235 ;
        RECT  0.305 -0.235 0.685 0.845 ;
        RECT  0.000 -0.235 0.305 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 3.685 3.360 4.155 ;
        RECT  1.970 2.780 2.350 4.155 ;
        RECT  0.685 3.685 1.970 4.155 ;
        RECT  0.305 2.595 0.685 4.155 ;
        RECT  0.000 3.685 0.305 4.155 ;
        END
    END VDD
END INVD3BWP7T

MACRO INVD4BWP7T
    CLASS CORE ;
    FOREIGN INVD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 0.495 2.895 1.375 ;
        RECT  2.610 2.175 2.840 3.350 ;
        RECT  2.410 2.175 2.610 2.525 ;
        RECT  2.410 1.025 2.555 1.375 ;
        RECT  1.510 1.025 2.410 2.525 ;
        RECT  1.390 1.025 1.510 1.375 ;
        RECT  1.330 2.175 1.510 2.525 ;
        RECT  1.045 0.490 1.390 1.375 ;
        RECT  1.100 2.175 1.330 3.350 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.605 1.280 1.945 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.665 -0.235 3.920 0.235 ;
        RECT  3.285 -0.235 3.665 1.190 ;
        RECT  2.160 -0.235 3.285 0.235 ;
        RECT  1.780 -0.235 2.160 0.795 ;
        RECT  0.685 -0.235 1.780 0.235 ;
        RECT  0.305 -0.235 0.685 0.845 ;
        RECT  0.000 -0.235 0.305 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.665 3.685 3.920 4.155 ;
        RECT  3.285 2.310 3.665 4.155 ;
        RECT  2.160 3.685 3.285 4.155 ;
        RECT  1.780 2.780 2.160 4.155 ;
        RECT  0.660 3.685 1.780 4.155 ;
        RECT  0.280 2.595 0.660 4.155 ;
        RECT  0.000 3.685 0.280 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.610 0.495 2.895 1.375 ;
        RECT  2.610 2.175 2.840 3.350 ;
        RECT  1.045 0.490 1.310 1.375 ;
        RECT  1.100 2.175 1.310 3.350 ;
    END
END INVD4BWP7T

MACRO INVD5BWP7T
    CLASS CORE ;
    FOREIGN INVD5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.6972 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.960 0.495 4.300 1.375 ;
        RECT  4.015 2.175 4.245 3.385 ;
        RECT  2.970 2.175 4.015 2.525 ;
        RECT  2.970 1.025 3.960 1.375 ;
        RECT  2.825 1.025 2.970 2.525 ;
        RECT  2.765 0.495 2.825 2.525 ;
        RECT  2.535 0.495 2.765 3.385 ;
        RECT  2.470 0.495 2.535 2.525 ;
        RECT  2.070 1.025 2.470 2.525 ;
        RECT  1.345 1.025 2.070 1.375 ;
        RECT  1.290 2.175 2.070 2.525 ;
        RECT  1.000 0.495 1.345 1.375 ;
        RECT  1.055 2.175 1.290 3.385 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 2.1330 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.605 1.820 1.945 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 -0.235 4.480 0.235 ;
        RECT  3.200 -0.235 3.580 0.795 ;
        RECT  2.100 -0.235 3.200 0.235 ;
        RECT  1.720 -0.235 2.100 0.795 ;
        RECT  0.620 -0.235 1.720 0.235 ;
        RECT  0.240 -0.235 0.620 0.945 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 3.685 4.480 4.155 ;
        RECT  3.200 2.780 3.580 4.155 ;
        RECT  2.100 3.685 3.200 4.155 ;
        RECT  1.720 2.780 2.100 4.155 ;
        RECT  0.620 3.685 1.720 4.155 ;
        RECT  0.240 2.595 0.620 4.155 ;
        RECT  0.000 3.685 0.240 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.960 0.495 4.300 1.375 ;
        RECT  4.015 2.175 4.245 3.385 ;
        RECT  3.170 2.175 4.015 2.525 ;
        RECT  3.170 1.025 3.960 1.375 ;
        RECT  1.345 1.025 1.870 1.375 ;
        RECT  1.290 2.175 1.870 2.525 ;
        RECT  1.000 0.495 1.345 1.375 ;
        RECT  1.055 2.175 1.290 3.385 ;
    END
END INVD5BWP7T

MACRO INVD6BWP7T
    CLASS CORE ;
    FOREIGN INVD6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.8394 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 0.495 4.120 1.375 ;
        RECT  3.835 2.175 4.065 3.410 ;
        RECT  2.970 2.175 3.835 2.525 ;
        RECT  2.970 1.025 3.780 1.375 ;
        RECT  2.690 1.025 2.970 2.525 ;
        RECT  2.625 0.495 2.690 2.525 ;
        RECT  2.395 0.495 2.625 3.410 ;
        RECT  2.340 0.495 2.395 2.525 ;
        RECT  2.070 1.025 2.340 2.525 ;
        RECT  1.250 1.025 2.070 1.375 ;
        RECT  1.185 2.175 2.070 2.525 ;
        RECT  0.900 0.490 1.250 1.375 ;
        RECT  0.955 2.175 1.185 3.410 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 2.5596 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.605 1.685 1.945 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.860 -0.235 5.040 0.235 ;
        RECT  4.480 -0.235 4.860 1.195 ;
        RECT  3.420 -0.235 4.480 0.235 ;
        RECT  3.040 -0.235 3.420 0.795 ;
        RECT  1.980 -0.235 3.040 0.235 ;
        RECT  1.600 -0.235 1.980 0.795 ;
        RECT  0.540 -0.235 1.600 0.235 ;
        RECT  0.160 -0.235 0.540 0.950 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.860 3.685 5.040 4.155 ;
        RECT  4.480 2.305 4.860 4.155 ;
        RECT  3.420 3.685 4.480 4.155 ;
        RECT  3.040 2.780 3.420 4.155 ;
        RECT  1.980 3.685 3.040 4.155 ;
        RECT  1.600 2.780 1.980 4.155 ;
        RECT  0.540 3.685 1.600 4.155 ;
        RECT  0.160 2.595 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 0.495 4.120 1.375 ;
        RECT  3.835 2.175 4.065 3.410 ;
        RECT  3.170 2.175 3.835 2.525 ;
        RECT  3.170 1.025 3.780 1.375 ;
        RECT  1.250 1.025 1.870 1.375 ;
        RECT  1.185 2.175 1.870 2.525 ;
        RECT  0.900 0.490 1.250 1.375 ;
        RECT  0.955 2.175 1.185 3.410 ;
    END
END INVD6BWP7T

MACRO INVD8BWP7T
    CLASS CORE ;
    FOREIGN INVD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.1192 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.375 0.490 5.720 1.400 ;
        RECT  5.430 2.150 5.660 3.435 ;
        RECT  4.200 2.150 5.430 2.550 ;
        RECT  4.255 1.000 5.375 1.400 ;
        RECT  4.090 0.490 4.255 1.400 ;
        RECT  4.090 2.150 4.200 3.435 ;
        RECT  3.970 0.490 4.090 3.435 ;
        RECT  3.910 0.490 3.970 2.550 ;
        RECT  3.190 1.000 3.910 2.550 ;
        RECT  2.795 1.000 3.190 1.400 ;
        RECT  2.740 2.150 3.190 2.550 ;
        RECT  2.455 0.490 2.795 1.400 ;
        RECT  2.510 2.150 2.740 3.435 ;
        RECT  1.280 2.150 2.510 2.550 ;
        RECT  1.335 1.000 2.455 1.400 ;
        RECT  0.995 0.490 1.335 1.400 ;
        RECT  1.050 2.150 1.280 3.435 ;
        END
    END ZN
    PIN I
        ANTENNAGATEAREA 3.4128 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.630 2.555 1.920 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END I
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 -0.235 6.720 0.235 ;
        RECT  6.105 -0.235 6.485 1.195 ;
        RECT  5.005 -0.235 6.105 0.235 ;
        RECT  4.625 -0.235 5.005 0.765 ;
        RECT  3.545 -0.235 4.625 0.235 ;
        RECT  3.165 -0.235 3.545 0.770 ;
        RECT  2.085 -0.235 3.165 0.235 ;
        RECT  1.705 -0.235 2.085 0.770 ;
        RECT  0.540 -0.235 1.705 0.235 ;
        RECT  0.160 -0.235 0.540 0.945 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 3.685 6.720 4.155 ;
        RECT  6.105 2.295 6.485 4.155 ;
        RECT  5.005 3.685 6.105 4.155 ;
        RECT  4.625 2.780 5.005 4.155 ;
        RECT  3.545 3.685 4.625 4.155 ;
        RECT  3.165 2.780 3.545 4.155 ;
        RECT  2.085 3.685 3.165 4.155 ;
        RECT  1.705 2.780 2.085 4.155 ;
        RECT  0.595 3.685 1.705 4.155 ;
        RECT  0.215 2.595 0.595 4.155 ;
        RECT  0.000 3.685 0.215 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.375 0.490 5.720 1.400 ;
        RECT  5.430 2.150 5.660 3.435 ;
        RECT  4.290 2.150 5.430 2.550 ;
        RECT  4.290 1.000 5.375 1.400 ;
        RECT  2.795 1.000 2.990 1.400 ;
        RECT  2.740 2.150 2.990 2.550 ;
        RECT  2.455 0.490 2.795 1.400 ;
        RECT  2.510 2.150 2.740 3.435 ;
        RECT  1.280 2.150 2.510 2.550 ;
        RECT  1.335 1.000 2.455 1.400 ;
        RECT  0.995 0.490 1.335 1.400 ;
        RECT  1.050 2.150 1.280 3.435 ;
    END
END INVD8BWP7T

MACRO IOA21D0BWP7T
    CLASS CORE ;
    FOREIGN IOA21D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6099 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 0.495 3.180 0.725 ;
        RECT  2.380 0.495 2.660 2.915 ;
        RECT  2.120 2.685 2.380 2.915 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.210 3.220 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.100 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.625 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.870 -0.235 3.360 0.235 ;
        RECT  1.490 -0.235 1.870 0.780 ;
        RECT  0.000 -0.235 1.490 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 3.685 3.360 4.155 ;
        RECT  2.895 2.650 3.125 4.155 ;
        RECT  1.640 3.685 2.895 4.155 ;
        RECT  1.255 3.455 1.640 4.155 ;
        RECT  0.550 3.685 1.255 4.155 ;
        RECT  0.140 3.455 0.550 4.155 ;
        RECT  0.000 3.685 0.140 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.920 1.135 2.085 1.365 ;
        RECT  0.910 2.595 1.085 2.825 ;
        RECT  0.910 0.535 0.920 1.365 ;
        RECT  0.680 0.535 0.910 2.825 ;
        RECT  0.185 0.535 0.680 0.765 ;
    END
END IOA21D0BWP7T

MACRO IOA21D1BWP7T
    CLASS CORE ;
    FOREIGN IOA21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2198 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 0.665 3.180 0.895 ;
        RECT  2.410 0.665 2.660 2.725 ;
        RECT  2.380 0.665 2.410 3.335 ;
        RECT  2.170 2.370 2.380 3.335 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.210 3.220 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.600 1.540 2.710 ;
        RECT  1.140 1.600 1.260 1.955 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.625 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.870 -0.235 3.360 0.235 ;
        RECT  1.490 -0.235 1.870 0.715 ;
        RECT  0.000 -0.235 1.490 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 3.685 3.360 4.155 ;
        RECT  2.895 2.505 3.125 4.155 ;
        RECT  1.640 3.685 2.895 4.155 ;
        RECT  1.255 3.455 1.640 4.155 ;
        RECT  0.550 3.685 1.255 4.155 ;
        RECT  0.140 3.455 0.550 4.155 ;
        RECT  0.000 3.685 0.140 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.820 1.135 2.055 1.965 ;
        RECT  0.920 1.135 1.820 1.365 ;
        RECT  0.910 2.420 1.030 2.760 ;
        RECT  0.910 0.515 0.920 1.365 ;
        RECT  0.680 0.515 0.910 2.760 ;
        RECT  0.185 0.515 0.680 0.745 ;
    END
END IOA21D1BWP7T

MACRO IOA21D2BWP7T
    CLASS CORE ;
    FOREIGN IOA21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.0196 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.835 2.470 4.065 3.420 ;
        RECT  3.780 2.470 3.835 2.710 ;
        RECT  3.500 0.925 3.780 2.710 ;
        RECT  3.060 0.925 3.500 1.155 ;
        RECT  2.625 2.470 3.500 2.710 ;
        RECT  2.395 2.470 2.625 3.420 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.660 3.240 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 1.680 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.790 -0.235 5.040 0.235 ;
        RECT  4.550 -0.235 4.790 1.275 ;
        RECT  1.910 -0.235 4.550 0.235 ;
        RECT  1.530 -0.235 1.910 0.790 ;
        RECT  0.000 -0.235 1.530 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.855 3.685 5.040 4.155 ;
        RECT  4.475 2.305 4.855 4.155 ;
        RECT  3.425 3.685 4.475 4.155 ;
        RECT  3.045 2.990 3.425 4.155 ;
        RECT  1.975 3.685 3.045 4.155 ;
        RECT  1.595 2.960 1.975 4.155 ;
        RECT  0.465 3.685 1.595 4.155 ;
        RECT  0.235 2.450 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.035 0.465 4.265 1.935 ;
        RECT  2.410 0.465 4.035 0.695 ;
        RECT  2.170 0.465 2.410 1.380 ;
        RECT  2.145 1.140 2.170 1.380 ;
        RECT  1.915 1.140 2.145 2.020 ;
        RECT  0.925 1.140 1.915 1.380 ;
        RECT  0.925 3.035 1.240 3.265 ;
        RECT  0.695 0.730 0.925 3.265 ;
        RECT  0.180 0.730 0.695 0.960 ;
    END
END IOA21D2BWP7T

MACRO IOA22D0BWP7T
    CLASS CORE ;
    FOREIGN IOA22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.8976 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 2.560 4.245 3.330 ;
        RECT  2.660 2.560 4.015 2.800 ;
        RECT  2.495 1.000 2.660 2.800 ;
        RECT  2.380 1.000 2.495 3.365 ;
        RECT  2.025 1.000 2.380 1.230 ;
        RECT  2.265 2.560 2.380 3.365 ;
        RECT  2.025 3.135 2.265 3.365 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.030 1.210 4.340 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 3.780 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.610 0.455 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.740 -0.235 4.480 0.235 ;
        RECT  3.360 -0.235 3.740 1.235 ;
        RECT  1.880 -0.235 3.360 0.235 ;
        RECT  1.510 -0.235 1.880 0.465 ;
        RECT  0.000 -0.235 1.510 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.030 3.685 4.480 4.155 ;
        RECT  2.800 3.040 3.030 4.155 ;
        RECT  1.665 3.685 2.800 4.155 ;
        RECT  1.320 3.450 1.665 4.155 ;
        RECT  0.525 3.685 1.320 4.155 ;
        RECT  0.185 3.450 0.525 4.155 ;
        RECT  0.000 3.685 0.185 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.010 1.655 2.135 1.885 ;
        RECT  1.780 1.655 2.010 2.845 ;
        RECT  0.935 2.615 1.780 2.845 ;
        RECT  0.705 0.935 0.935 2.845 ;
        RECT  0.465 0.935 0.705 1.175 ;
        RECT  0.235 0.520 0.465 1.175 ;
    END
END IOA22D0BWP7T

MACRO IOA22D1BWP7T
    CLASS CORE ;
    FOREIGN IOA22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8774 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 2.425 4.690 3.275 ;
        RECT  2.660 2.425 4.450 2.665 ;
        RECT  2.645 0.485 2.660 2.665 ;
        RECT  2.380 0.485 2.645 3.325 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.620 4.900 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.675 3.800 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2466 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.620 0.465 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2466 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 1.210 1.540 2.190 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 -0.235 5.040 0.235 ;
        RECT  3.780 -0.235 4.160 0.845 ;
        RECT  1.930 -0.235 3.780 0.235 ;
        RECT  1.575 -0.235 1.930 0.470 ;
        RECT  0.000 -0.235 1.575 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 3.685 5.040 4.155 ;
        RECT  3.060 2.935 3.440 4.155 ;
        RECT  2.005 3.685 3.060 4.155 ;
        RECT  1.655 3.420 2.005 4.155 ;
        RECT  0.540 3.685 1.655 4.155 ;
        RECT  0.160 3.015 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.575 0.495 4.805 1.355 ;
        RECT  3.365 1.115 4.575 1.355 ;
        RECT  3.135 0.495 3.365 1.355 ;
        RECT  1.865 0.725 2.095 3.175 ;
        RECT  0.180 0.725 1.865 0.955 ;
        RECT  0.900 2.945 1.865 3.175 ;
    END
END IOA22D1BWP7T

MACRO IOA22D2BWP7T
    CLASS CORE ;
    FOREIGN IOA22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.925 4.340 2.710 ;
        RECT  3.515 0.925 4.060 1.155 ;
        RECT  3.910 2.415 4.060 2.710 ;
        RECT  3.680 2.415 3.910 3.385 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.710 1.540 6.020 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 2.000 3.220 2.710 ;
        RECT  2.660 2.000 2.940 2.230 ;
        RECT  2.380 1.615 2.660 2.230 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.660 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 -0.235 6.160 0.235 ;
        RECT  5.695 -0.235 5.925 1.230 ;
        RECT  2.800 -0.235 5.695 0.235 ;
        RECT  2.460 -0.235 2.800 0.465 ;
        RECT  0.520 -0.235 2.460 0.235 ;
        RECT  0.180 -0.235 0.520 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.700 3.685 6.160 4.155 ;
        RECT  4.320 3.080 4.700 4.155 ;
        RECT  3.190 3.685 4.320 4.155 ;
        RECT  2.955 3.150 3.190 4.155 ;
        RECT  1.980 3.685 2.955 4.155 ;
        RECT  1.600 3.125 1.980 4.155 ;
        RECT  0.000 3.685 1.600 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.465 2.940 5.980 3.170 ;
        RECT  5.235 0.980 5.465 3.170 ;
        RECT  5.065 0.980 5.235 1.210 ;
        RECT  4.835 0.465 5.065 1.210 ;
        RECT  3.260 0.465 4.835 0.695 ;
        RECT  3.180 1.540 3.755 1.770 ;
        RECT  3.030 0.465 3.260 0.925 ;
        RECT  2.950 1.155 3.180 1.770 ;
        RECT  2.065 0.695 3.030 0.925 ;
        RECT  1.440 1.155 2.950 1.385 ;
        RECT  2.405 2.475 2.635 2.875 ;
        RECT  1.185 2.645 2.405 2.875 ;
        RECT  1.835 0.465 2.065 0.925 ;
        RECT  0.980 0.465 1.835 0.695 ;
        RECT  1.210 0.965 1.440 1.385 ;
        RECT  1.020 1.155 1.210 1.385 ;
        RECT  0.955 2.645 1.185 3.455 ;
        RECT  0.780 1.155 1.020 2.400 ;
        RECT  0.750 0.465 0.980 0.925 ;
        RECT  0.465 2.170 0.780 2.400 ;
        RECT  0.520 0.695 0.750 0.925 ;
        RECT  0.290 0.695 0.520 1.940 ;
        RECT  0.230 2.170 0.465 3.380 ;
    END
END IOA22D2BWP7T

MACRO LHCND1BWP7T
    CLASS CORE ;
    FOREIGN LHCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.0426 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.020 9.380 2.530 ;
        RECT  8.680 1.020 9.100 1.250 ;
        RECT  8.680 2.300 9.100 2.530 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.175 0.495 10.500 3.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.650 3.235 1.790 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.3393 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.650 2.660 1.790 ;
        RECT  2.335 1.450 2.380 1.790 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.755 -0.235 10.640 0.235 ;
        RECT  9.375 -0.235 9.755 0.775 ;
        RECT  7.560 -0.235 9.375 0.235 ;
        RECT  7.220 -0.235 7.560 0.570 ;
        RECT  6.450 -0.235 7.220 0.235 ;
        RECT  6.220 -0.235 6.450 1.215 ;
        RECT  2.150 -0.235 6.220 0.235 ;
        RECT  5.935 0.985 6.220 1.215 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.740 3.685 10.640 4.155 ;
        RECT  9.400 3.220 9.740 4.155 ;
        RECT  7.685 3.685 9.400 4.155 ;
        RECT  7.345 3.245 7.685 4.155 ;
        RECT  6.370 3.685 7.345 4.155 ;
        RECT  6.140 3.160 6.370 4.155 ;
        RECT  3.245 3.685 6.140 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.695 1.660 9.925 2.990 ;
        RECT  8.365 2.760 9.695 2.990 ;
        RECT  8.135 0.465 8.365 3.440 ;
        RECT  7.980 0.465 8.135 0.695 ;
        RECT  7.090 1.700 7.855 2.040 ;
        RECT  6.860 0.965 7.090 2.930 ;
        RECT  6.735 0.965 6.860 1.305 ;
        RECT  5.850 2.700 6.860 2.930 ;
        RECT  5.390 1.755 6.515 1.985 ;
        RECT  5.620 2.700 5.850 3.455 ;
        RECT  5.160 0.985 5.390 3.455 ;
        RECT  4.220 0.985 5.160 1.215 ;
        RECT  3.785 3.225 5.160 3.455 ;
        RECT  4.700 1.505 4.930 2.990 ;
        RECT  3.775 1.505 4.700 1.735 ;
        RECT  4.040 2.120 4.270 2.710 ;
        RECT  2.325 2.480 4.040 2.710 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  3.545 1.505 3.775 2.250 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  1.840 2.020 3.545 2.250 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 1.020 1.840 2.535 ;
        RECT  1.500 1.020 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LHCND1BWP7T

MACRO LHCND2BWP7T
    CLASS CORE ;
    FOREIGN LHCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.2848 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.640 0.495 9.980 2.530 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.365 1.210 11.620 2.450 ;
        RECT  11.340 0.495 11.365 3.275 ;
        RECT  11.135 0.495 11.340 1.440 ;
        RECT  11.135 2.220 11.340 3.275 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.650 3.235 1.790 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.2952 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.650 2.660 1.790 ;
        RECT  2.335 1.450 2.380 1.790 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.085 -0.235 12.320 0.235 ;
        RECT  11.855 -0.235 12.085 1.260 ;
        RECT  10.725 -0.235 11.855 0.235 ;
        RECT  10.345 -0.235 10.725 0.910 ;
        RECT  9.125 -0.235 10.345 0.235 ;
        RECT  8.895 -0.235 9.125 1.235 ;
        RECT  7.720 -0.235 8.895 0.235 ;
        RECT  7.380 -0.235 7.720 1.165 ;
        RECT  6.450 -0.235 7.380 0.235 ;
        RECT  6.220 -0.235 6.450 1.215 ;
        RECT  2.150 -0.235 6.220 0.235 ;
        RECT  5.935 0.985 6.220 1.215 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.085 3.685 12.320 4.155 ;
        RECT  11.855 2.250 12.085 4.155 ;
        RECT  10.720 3.685 11.855 4.155 ;
        RECT  10.340 3.250 10.720 4.155 ;
        RECT  9.260 3.685 10.340 4.155 ;
        RECT  8.920 3.250 9.260 4.155 ;
        RECT  7.840 3.685 8.920 4.155 ;
        RECT  7.500 2.305 7.840 4.155 ;
        RECT  6.365 3.685 7.500 4.155 ;
        RECT  6.135 3.160 6.365 4.155 ;
        RECT  3.245 3.685 6.135 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.655 1.620 10.885 3.020 ;
        RECT  8.505 2.790 10.655 3.020 ;
        RECT  8.275 0.495 8.505 3.125 ;
        RECT  8.190 0.495 8.275 1.305 ;
        RECT  7.090 1.660 8.015 2.000 ;
        RECT  6.855 0.495 7.090 3.085 ;
        RECT  6.735 0.495 6.855 1.305 ;
        RECT  5.845 2.700 6.855 2.930 ;
        RECT  5.385 1.755 6.515 1.985 ;
        RECT  5.615 2.700 5.845 3.455 ;
        RECT  5.155 0.985 5.385 3.455 ;
        RECT  4.220 0.985 5.155 1.215 ;
        RECT  3.785 3.225 5.155 3.455 ;
        RECT  4.695 1.515 4.925 2.990 ;
        RECT  4.040 1.515 4.695 1.745 ;
        RECT  4.040 2.120 4.270 2.710 ;
        RECT  3.775 1.505 4.040 1.745 ;
        RECT  2.325 2.480 4.040 2.710 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  3.545 1.505 3.775 2.250 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  1.840 2.020 3.545 2.250 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 1.020 1.840 2.535 ;
        RECT  1.500 1.020 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LHCND2BWP7T

MACRO LHCNQD1BWP7T
    CLASS CORE ;
    FOREIGN LHCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.615 0.495 9.940 3.300 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.650 3.235 1.790 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.3393 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.650 2.660 1.790 ;
        RECT  2.335 1.450 2.380 1.790 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.195 -0.235 10.080 0.235 ;
        RECT  8.815 -0.235 9.195 1.140 ;
        RECT  7.760 -0.235 8.815 0.235 ;
        RECT  7.420 -0.235 7.760 1.140 ;
        RECT  6.450 -0.235 7.420 0.235 ;
        RECT  6.220 -0.235 6.450 1.215 ;
        RECT  2.150 -0.235 6.220 0.235 ;
        RECT  5.935 0.985 6.220 1.215 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.180 3.685 10.080 4.155 ;
        RECT  8.840 2.310 9.180 4.155 ;
        RECT  7.745 3.685 8.840 4.155 ;
        RECT  7.405 3.245 7.745 4.155 ;
        RECT  6.370 3.685 7.405 4.155 ;
        RECT  6.140 3.160 6.370 4.155 ;
        RECT  3.245 3.685 6.140 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.425 1.660 9.365 2.000 ;
        RECT  8.195 0.465 8.425 3.440 ;
        RECT  7.090 1.700 7.915 2.040 ;
        RECT  6.860 0.965 7.090 2.930 ;
        RECT  6.735 0.965 6.860 1.305 ;
        RECT  5.850 2.700 6.860 2.930 ;
        RECT  5.390 1.755 6.515 1.985 ;
        RECT  5.620 2.700 5.850 3.455 ;
        RECT  5.160 0.985 5.390 3.455 ;
        RECT  4.220 0.985 5.160 1.215 ;
        RECT  3.785 3.225 5.160 3.455 ;
        RECT  4.700 1.515 4.930 2.990 ;
        RECT  4.040 1.515 4.700 1.745 ;
        RECT  4.040 2.120 4.270 2.710 ;
        RECT  3.775 1.505 4.040 1.745 ;
        RECT  2.325 2.480 4.040 2.710 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  3.545 1.505 3.775 2.250 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  1.840 2.020 3.545 2.250 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 1.020 1.840 2.535 ;
        RECT  1.500 1.020 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LHCNQD1BWP7T

MACRO LHCNQD2BWP7T
    CLASS CORE ;
    FOREIGN LHCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.125 1.210 9.380 2.450 ;
        RECT  9.100 0.495 9.125 3.275 ;
        RECT  8.895 0.495 9.100 1.440 ;
        RECT  8.895 2.220 9.100 3.275 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.650 3.235 1.790 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.2952 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.650 2.660 1.790 ;
        RECT  2.335 1.450 2.380 1.790 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 -0.235 10.080 0.235 ;
        RECT  9.615 -0.235 9.845 1.260 ;
        RECT  8.485 -0.235 9.615 0.235 ;
        RECT  8.105 -0.235 8.485 0.670 ;
        RECT  6.450 -0.235 8.105 0.235 ;
        RECT  6.220 -0.235 6.450 1.215 ;
        RECT  2.150 -0.235 6.220 0.235 ;
        RECT  5.935 0.985 6.220 1.215 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 3.685 10.080 4.155 ;
        RECT  9.615 2.250 9.845 4.155 ;
        RECT  8.480 3.685 9.615 4.155 ;
        RECT  8.100 3.250 8.480 4.155 ;
        RECT  6.365 3.685 8.100 4.155 ;
        RECT  6.135 3.160 6.365 4.155 ;
        RECT  3.245 3.685 6.135 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.415 1.075 8.645 3.000 ;
        RECT  7.685 1.075 8.415 1.305 ;
        RECT  7.685 2.770 8.415 3.000 ;
        RECT  7.090 1.660 7.915 2.000 ;
        RECT  7.455 0.495 7.685 1.305 ;
        RECT  7.455 2.770 7.685 3.440 ;
        RECT  6.855 0.495 7.090 2.930 ;
        RECT  6.735 0.495 6.855 1.305 ;
        RECT  5.845 2.700 6.855 2.930 ;
        RECT  5.385 1.755 6.515 1.985 ;
        RECT  5.615 2.700 5.845 3.455 ;
        RECT  5.155 0.985 5.385 3.455 ;
        RECT  4.220 0.985 5.155 1.215 ;
        RECT  3.785 3.225 5.155 3.455 ;
        RECT  4.695 1.515 4.925 2.990 ;
        RECT  4.040 1.515 4.695 1.745 ;
        RECT  4.040 2.120 4.270 2.710 ;
        RECT  3.775 1.505 4.040 1.745 ;
        RECT  2.325 2.480 4.040 2.710 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  3.545 1.505 3.775 2.250 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  1.840 2.020 3.545 2.250 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 1.020 1.840 2.535 ;
        RECT  1.500 1.020 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LHCNQD2BWP7T

MACRO LHD1BWP7T
    CLASS CORE ;
    FOREIGN LHD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.935 0.495 8.260 3.300 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.0040 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.580 0.495 6.730 1.305 ;
        RECT  6.580 2.415 6.700 2.645 ;
        RECT  6.300 0.495 6.580 2.645 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.475 -0.235 8.400 0.235 ;
        RECT  7.095 -0.235 7.475 0.940 ;
        RECT  5.200 -0.235 7.095 0.235 ;
        RECT  4.820 -0.235 5.200 0.670 ;
        RECT  2.420 -0.235 4.820 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.460 3.685 8.400 4.155 ;
        RECT  7.120 3.455 7.460 4.155 ;
        RECT  5.290 3.685 7.120 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.455 1.660 7.685 3.190 ;
        RECT  6.010 2.960 7.455 3.190 ;
        RECT  5.850 1.295 6.010 3.440 ;
        RECT  5.780 0.965 5.850 3.440 ;
        RECT  5.620 0.965 5.780 1.525 ;
        RECT  4.465 1.295 5.620 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.275 3.775 2.720 ;
        RECT  3.260 1.275 3.545 1.505 ;
        RECT  3.220 1.900 3.315 2.240 ;
        RECT  3.030 0.930 3.260 1.505 ;
        RECT  2.990 1.900 3.220 3.210 ;
        RECT  2.080 0.930 3.030 1.160 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  1.850 0.930 2.080 2.720 ;
        RECT  1.500 0.930 1.850 1.160 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LHD1BWP7T

MACRO LHD2BWP7T
    CLASS CORE ;
    FOREIGN LHD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.155 9.380 2.485 ;
        RECT  8.860 1.155 9.100 1.385 ;
        RECT  8.860 2.255 9.100 2.485 ;
        RECT  8.630 0.485 8.860 1.385 ;
        RECT  8.630 2.255 8.860 3.205 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.420 1.075 7.700 2.530 ;
        RECT  7.190 0.495 7.420 1.305 ;
        RECT  7.135 2.255 7.420 2.530 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 -0.235 10.080 0.235 ;
        RECT  9.615 -0.235 9.845 1.250 ;
        RECT  8.225 -0.235 9.615 0.235 ;
        RECT  7.845 -0.235 8.225 0.820 ;
        RECT  6.715 -0.235 7.845 0.235 ;
        RECT  6.375 -0.235 6.715 1.225 ;
        RECT  5.200 -0.235 6.375 0.235 ;
        RECT  4.820 -0.235 5.200 0.670 ;
        RECT  2.420 -0.235 4.820 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 3.685 10.080 4.155 ;
        RECT  9.615 2.255 9.845 4.155 ;
        RECT  8.265 3.685 9.615 4.155 ;
        RECT  7.805 3.250 8.265 4.155 ;
        RECT  6.765 3.685 7.805 4.155 ;
        RECT  6.305 3.250 6.765 4.155 ;
        RECT  5.290 3.685 6.305 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.320 1.715 8.715 1.945 ;
        RECT  8.040 1.715 8.320 3.020 ;
        RECT  6.010 2.790 8.040 3.020 ;
        RECT  5.960 1.295 6.010 3.020 ;
        RECT  5.780 0.495 5.960 3.020 ;
        RECT  5.730 0.495 5.780 1.525 ;
        RECT  4.465 1.295 5.730 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.275 3.775 2.720 ;
        RECT  3.260 1.275 3.545 1.505 ;
        RECT  3.220 1.900 3.315 2.240 ;
        RECT  3.030 0.930 3.260 1.505 ;
        RECT  2.990 1.900 3.220 3.210 ;
        RECT  2.080 0.930 3.030 1.160 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  1.850 0.930 2.080 2.720 ;
        RECT  1.500 0.930 1.850 1.160 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LHD2BWP7T

MACRO LHQD1BWP7T
    CLASS CORE ;
    FOREIGN LHQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.180 7.140 2.480 ;
        RECT  6.730 1.180 6.860 1.410 ;
        RECT  6.730 2.250 6.860 2.480 ;
        RECT  6.500 0.495 6.730 1.410 ;
        RECT  6.500 2.250 6.730 3.200 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.605 -0.235 7.840 0.235 ;
        RECT  7.375 -0.235 7.605 1.235 ;
        RECT  7.225 -0.235 7.375 0.420 ;
        RECT  5.200 -0.235 7.225 0.235 ;
        RECT  4.820 -0.235 5.200 0.670 ;
        RECT  2.420 -0.235 4.820 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.600 3.685 7.840 4.155 ;
        RECT  7.370 2.245 7.600 4.155 ;
        RECT  5.290 3.685 7.370 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.780 0.495 6.010 3.200 ;
        RECT  4.465 1.295 5.780 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.275 3.775 2.720 ;
        RECT  3.260 1.275 3.545 1.505 ;
        RECT  3.220 1.900 3.315 2.240 ;
        RECT  3.030 0.930 3.260 1.505 ;
        RECT  2.990 1.900 3.220 3.210 ;
        RECT  2.080 0.930 3.030 1.160 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  1.850 0.930 2.080 2.720 ;
        RECT  1.500 0.930 1.850 1.160 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LHQD1BWP7T

MACRO LHQD2BWP7T
    CLASS CORE ;
    FOREIGN LHQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.445 1.180 7.700 2.480 ;
        RECT  7.420 0.495 7.445 3.200 ;
        RECT  7.215 0.495 7.420 1.410 ;
        RECT  7.215 2.250 7.420 3.200 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.165 -0.235 8.400 0.235 ;
        RECT  7.935 -0.235 8.165 1.250 ;
        RECT  6.795 -0.235 7.935 0.235 ;
        RECT  6.415 -0.235 6.795 1.205 ;
        RECT  5.200 -0.235 6.415 0.235 ;
        RECT  4.820 -0.235 5.200 0.670 ;
        RECT  2.420 -0.235 4.820 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.165 3.685 8.400 4.155 ;
        RECT  7.935 2.245 8.165 4.155 ;
        RECT  6.795 3.685 7.935 4.155 ;
        RECT  6.415 2.310 6.795 4.155 ;
        RECT  5.290 3.685 6.415 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.780 0.495 6.010 3.200 ;
        RECT  4.465 1.295 5.780 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.275 3.775 2.720 ;
        RECT  3.260 1.275 3.545 1.505 ;
        RECT  3.220 1.900 3.315 2.240 ;
        RECT  3.030 0.930 3.260 1.505 ;
        RECT  2.990 1.900 3.220 3.210 ;
        RECT  2.080 0.930 3.030 1.160 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  1.850 0.930 2.080 2.720 ;
        RECT  1.500 0.930 1.850 1.160 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LHQD2BWP7T

MACRO LHSND1BWP7T
    CLASS CORE ;
    FOREIGN LHSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3087 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.615 0.495 9.940 3.185 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.075 8.820 2.535 ;
        RECT  8.405 1.075 8.540 1.305 ;
        RECT  8.120 2.305 8.540 2.535 ;
        RECT  8.175 0.485 8.405 1.305 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 1.210 2.680 2.150 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.240 -0.235 10.080 0.235 ;
        RECT  8.780 -0.235 9.240 0.845 ;
        RECT  6.985 -0.235 8.780 0.235 ;
        RECT  6.755 -0.235 6.985 0.840 ;
        RECT  5.140 -0.235 6.755 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.250 3.685 10.080 4.155 ;
        RECT  8.790 3.250 9.250 4.155 ;
        RECT  6.800 3.685 8.790 4.155 ;
        RECT  6.455 3.445 6.800 4.155 ;
        RECT  2.545 3.685 6.455 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.135 1.660 9.365 3.020 ;
        RECT  7.035 2.790 9.135 3.020 ;
        RECT  7.710 1.590 8.310 1.935 ;
        RECT  7.430 0.500 7.710 2.560 ;
        RECT  7.290 2.330 7.430 2.560 ;
        RECT  6.805 1.160 7.035 3.020 ;
        RECT  6.480 1.160 6.805 1.390 ;
        RECT  5.980 2.790 6.805 3.020 ;
        RECT  6.250 0.605 6.480 1.390 ;
        RECT  5.990 0.605 6.250 0.835 ;
        RECT  5.750 2.790 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.935 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.655 2.705 4.875 2.935 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.290 1.070 3.760 1.300 ;
        RECT  3.315 1.685 3.530 2.400 ;
        RECT  3.300 1.685 3.315 3.170 ;
        RECT  3.075 2.170 3.300 3.170 ;
        RECT  3.060 0.750 3.290 1.300 ;
        RECT  1.455 2.940 3.075 3.170 ;
        RECT  2.060 0.750 3.060 0.980 ;
        RECT  1.830 0.750 2.060 2.710 ;
        RECT  1.760 0.750 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LHSND1BWP7T

MACRO LHSND2BWP7T
    CLASS CORE ;
    FOREIGN LHSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.2988 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.780 1.210 11.060 2.450 ;
        RECT  10.685 1.210 10.780 1.440 ;
        RECT  10.685 2.220 10.780 2.450 ;
        RECT  10.455 0.495 10.685 1.440 ;
        RECT  10.455 2.220 10.685 3.275 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.4898 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.870 0.495 9.100 1.400 ;
        RECT  8.820 2.300 9.075 2.530 ;
        RECT  8.820 1.165 8.870 1.400 ;
        RECT  8.540 1.165 8.820 2.530 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.3321 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 1.210 2.680 2.150 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.525 -0.235 11.760 0.235 ;
        RECT  11.295 -0.235 11.525 1.260 ;
        RECT  10.030 -0.235 11.295 0.235 ;
        RECT  9.650 -0.235 10.030 0.910 ;
        RECT  8.210 -0.235 9.650 0.235 ;
        RECT  7.980 -0.235 8.210 1.235 ;
        RECT  5.140 -0.235 7.980 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.520 3.685 11.760 4.155 ;
        RECT  11.290 2.250 11.520 4.155 ;
        RECT  9.925 3.685 11.290 4.155 ;
        RECT  9.545 3.250 9.925 4.155 ;
        RECT  8.355 3.685 9.545 4.155 ;
        RECT  8.015 3.250 8.355 4.155 ;
        RECT  6.880 3.685 8.015 4.155 ;
        RECT  6.485 3.455 6.880 4.155 ;
        RECT  2.545 3.685 6.485 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.975 1.620 10.205 3.020 ;
        RECT  7.060 2.790 9.975 3.020 ;
        RECT  7.710 1.655 8.290 2.030 ;
        RECT  7.430 0.585 7.710 2.530 ;
        RECT  7.075 0.585 7.430 0.815 ;
        RECT  7.290 2.300 7.430 2.530 ;
        RECT  6.830 1.110 7.060 3.020 ;
        RECT  6.670 1.110 6.830 1.340 ;
        RECT  5.980 2.790 6.830 3.020 ;
        RECT  6.440 0.605 6.670 1.340 ;
        RECT  5.990 0.605 6.440 0.835 ;
        RECT  5.750 2.790 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.935 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.655 2.705 4.875 2.935 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.285 1.070 3.760 1.300 ;
        RECT  3.315 1.625 3.530 2.400 ;
        RECT  3.300 1.625 3.315 3.170 ;
        RECT  3.075 2.170 3.300 3.170 ;
        RECT  3.055 0.750 3.285 1.300 ;
        RECT  1.455 2.940 3.075 3.170 ;
        RECT  2.060 0.750 3.055 0.980 ;
        RECT  1.830 0.750 2.060 2.710 ;
        RECT  1.760 0.750 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LHSND2BWP7T

MACRO LHSNQD1BWP7T
    CLASS CORE ;
    FOREIGN LHSNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3033 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.5168 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.055 0.485 9.385 3.195 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2700 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 1.210 2.680 2.150 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.520 -0.235 9.520 0.235 ;
        RECT  8.060 -0.235 8.520 1.140 ;
        RECT  6.985 -0.235 8.060 0.235 ;
        RECT  6.755 -0.235 6.985 0.840 ;
        RECT  5.140 -0.235 6.755 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.530 3.685 9.520 4.155 ;
        RECT  8.070 2.310 8.530 4.155 ;
        RECT  6.800 3.685 8.070 4.155 ;
        RECT  6.455 3.445 6.800 4.155 ;
        RECT  2.545 3.685 6.455 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.710 1.590 8.645 1.935 ;
        RECT  7.430 0.500 7.710 2.560 ;
        RECT  7.290 2.330 7.430 2.560 ;
        RECT  6.805 1.160 7.035 3.020 ;
        RECT  6.480 1.160 6.805 1.390 ;
        RECT  5.980 2.790 6.805 3.020 ;
        RECT  6.250 0.605 6.480 1.390 ;
        RECT  5.990 0.605 6.250 0.835 ;
        RECT  5.750 2.790 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.935 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.655 2.705 4.875 2.935 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.285 1.070 3.760 1.300 ;
        RECT  3.315 1.685 3.530 2.400 ;
        RECT  3.300 1.685 3.315 3.170 ;
        RECT  3.075 2.170 3.300 3.170 ;
        RECT  3.055 0.750 3.285 1.300 ;
        RECT  1.455 2.940 3.075 3.170 ;
        RECT  2.060 0.750 3.055 0.980 ;
        RECT  1.830 0.750 2.060 2.710 ;
        RECT  1.760 0.750 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LHSNQD1BWP7T

MACRO LHSNQD2BWP7T
    CLASS CORE ;
    FOREIGN LHSNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.2988 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.4098 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.870 0.495 9.100 1.400 ;
        RECT  8.820 2.245 9.025 3.200 ;
        RECT  8.820 1.165 8.870 1.400 ;
        RECT  8.790 1.165 8.820 3.200 ;
        RECT  8.540 1.165 8.790 2.530 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2700 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 1.210 2.680 2.150 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.900 -0.235 10.080 0.235 ;
        RECT  9.560 -0.235 9.900 1.180 ;
        RECT  8.210 -0.235 9.560 0.235 ;
        RECT  7.980 -0.235 8.210 1.235 ;
        RECT  5.140 -0.235 7.980 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.920 3.685 10.080 4.155 ;
        RECT  9.540 2.310 9.920 4.155 ;
        RECT  8.300 3.685 9.540 4.155 ;
        RECT  8.070 2.255 8.300 4.155 ;
        RECT  6.880 3.685 8.070 4.155 ;
        RECT  6.485 3.455 6.880 4.155 ;
        RECT  2.545 3.685 6.485 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.710 1.655 8.290 2.000 ;
        RECT  7.430 0.585 7.710 2.530 ;
        RECT  7.075 0.585 7.430 0.815 ;
        RECT  7.290 2.300 7.430 2.530 ;
        RECT  6.830 1.110 7.060 3.020 ;
        RECT  6.670 1.110 6.830 1.340 ;
        RECT  5.980 2.790 6.830 3.020 ;
        RECT  6.440 0.605 6.670 1.340 ;
        RECT  5.990 0.605 6.440 0.835 ;
        RECT  5.750 2.790 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.970 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.655 2.740 4.875 2.970 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.285 1.070 3.760 1.300 ;
        RECT  3.315 1.685 3.530 2.400 ;
        RECT  3.300 1.685 3.315 3.170 ;
        RECT  3.075 2.170 3.300 3.170 ;
        RECT  3.055 0.750 3.285 1.300 ;
        RECT  1.455 2.940 3.075 3.170 ;
        RECT  2.060 0.750 3.055 0.980 ;
        RECT  1.830 0.750 2.060 2.710 ;
        RECT  1.760 0.750 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LHSNQD2BWP7T

MACRO LNCND1BWP7T
    CLASS CORE ;
    FOREIGN LNCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.0426 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.020 9.380 2.530 ;
        RECT  8.680 1.020 9.100 1.250 ;
        RECT  8.680 2.300 9.100 2.530 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.175 0.495 10.500 3.300 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3042 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.235 2.150 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.330 1.485 2.380 1.825 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.755 -0.235 10.640 0.235 ;
        RECT  9.375 -0.235 9.755 0.775 ;
        RECT  7.560 -0.235 9.375 0.235 ;
        RECT  7.220 -0.235 7.560 0.570 ;
        RECT  6.450 -0.235 7.220 0.235 ;
        RECT  6.220 -0.235 6.450 1.215 ;
        RECT  2.150 -0.235 6.220 0.235 ;
        RECT  5.935 0.985 6.220 1.215 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.740 3.685 10.640 4.155 ;
        RECT  9.400 3.220 9.740 4.155 ;
        RECT  7.685 3.685 9.400 4.155 ;
        RECT  7.345 3.245 7.685 4.155 ;
        RECT  6.370 3.685 7.345 4.155 ;
        RECT  6.140 3.160 6.370 4.155 ;
        RECT  3.245 3.685 6.140 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.695 1.660 9.925 2.990 ;
        RECT  8.365 2.760 9.695 2.990 ;
        RECT  8.135 0.465 8.365 3.440 ;
        RECT  7.980 0.465 8.135 0.695 ;
        RECT  7.090 1.700 7.855 2.040 ;
        RECT  6.860 0.965 7.090 2.930 ;
        RECT  6.735 0.965 6.860 1.305 ;
        RECT  5.850 2.700 6.860 2.930 ;
        RECT  6.230 1.700 6.460 2.250 ;
        RECT  5.390 2.020 6.230 2.250 ;
        RECT  5.620 2.700 5.850 3.455 ;
        RECT  5.160 2.020 5.390 3.455 ;
        RECT  4.365 2.020 5.160 2.250 ;
        RECT  3.785 3.225 5.160 3.455 ;
        RECT  4.705 0.525 4.935 1.790 ;
        RECT  4.700 2.480 4.930 2.990 ;
        RECT  3.820 0.525 4.705 0.755 ;
        RECT  4.595 1.450 4.705 1.790 ;
        RECT  3.905 2.480 4.700 2.710 ;
        RECT  4.365 0.985 4.475 1.215 ;
        RECT  4.135 0.985 4.365 2.250 ;
        RECT  3.675 1.485 3.905 2.710 ;
        RECT  3.590 0.525 3.820 0.925 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  2.325 2.480 3.675 2.710 ;
        RECT  1.840 0.695 3.590 0.925 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 0.695 1.840 2.535 ;
        RECT  1.500 0.695 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LNCND1BWP7T

MACRO LNCND2BWP7T
    CLASS CORE ;
    FOREIGN LNCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.2848 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.640 0.495 9.980 2.530 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.365 1.210 11.620 2.450 ;
        RECT  11.340 0.495 11.365 3.275 ;
        RECT  11.135 0.495 11.340 1.440 ;
        RECT  11.135 2.220 11.340 3.275 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3042 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.235 2.150 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.330 1.485 2.380 1.825 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.085 -0.235 12.320 0.235 ;
        RECT  11.855 -0.235 12.085 1.260 ;
        RECT  10.725 -0.235 11.855 0.235 ;
        RECT  10.345 -0.235 10.725 0.910 ;
        RECT  9.125 -0.235 10.345 0.235 ;
        RECT  8.895 -0.235 9.125 1.235 ;
        RECT  7.740 -0.235 8.895 0.235 ;
        RECT  7.400 -0.235 7.740 1.140 ;
        RECT  6.285 -0.235 7.400 0.235 ;
        RECT  5.935 -0.235 6.285 1.215 ;
        RECT  2.150 -0.235 5.935 0.235 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.085 3.685 12.320 4.155 ;
        RECT  11.855 2.250 12.085 4.155 ;
        RECT  10.720 3.685 11.855 4.155 ;
        RECT  10.340 3.250 10.720 4.155 ;
        RECT  9.260 3.685 10.340 4.155 ;
        RECT  8.920 3.250 9.260 4.155 ;
        RECT  7.840 3.685 8.920 4.155 ;
        RECT  7.500 2.305 7.840 4.155 ;
        RECT  6.420 3.685 7.500 4.155 ;
        RECT  6.080 3.245 6.420 4.155 ;
        RECT  3.245 3.685 6.080 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.655 1.620 10.885 3.020 ;
        RECT  8.505 2.790 10.655 3.020 ;
        RECT  8.275 0.495 8.505 3.095 ;
        RECT  8.120 0.495 8.275 1.305 ;
        RECT  7.085 1.660 7.995 2.000 ;
        RECT  6.855 0.495 7.085 3.095 ;
        RECT  6.735 0.495 6.855 1.305 ;
        RECT  5.845 2.785 6.855 3.015 ;
        RECT  6.230 1.700 6.460 2.250 ;
        RECT  5.385 2.020 6.230 2.250 ;
        RECT  5.615 2.785 5.845 3.455 ;
        RECT  5.155 2.020 5.385 3.455 ;
        RECT  4.365 2.020 5.155 2.250 ;
        RECT  3.785 3.225 5.155 3.455 ;
        RECT  4.705 0.525 4.935 1.790 ;
        RECT  4.695 2.480 4.925 2.990 ;
        RECT  3.820 0.525 4.705 0.755 ;
        RECT  4.595 1.450 4.705 1.790 ;
        RECT  3.905 2.480 4.695 2.710 ;
        RECT  4.365 0.985 4.475 1.215 ;
        RECT  4.135 0.985 4.365 2.250 ;
        RECT  3.675 1.485 3.905 2.710 ;
        RECT  3.590 0.525 3.820 0.925 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  2.325 2.480 3.675 2.710 ;
        RECT  1.840 0.695 3.590 0.925 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 0.695 1.840 2.535 ;
        RECT  1.500 0.695 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LNCND2BWP7T

MACRO LNCNQD1BWP7T
    CLASS CORE ;
    FOREIGN LNCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.055 0.495 9.380 3.300 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3042 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.235 2.150 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.330 1.485 2.380 1.825 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.635 -0.235 9.520 0.235 ;
        RECT  8.255 -0.235 8.635 1.140 ;
        RECT  6.370 -0.235 8.255 0.235 ;
        RECT  6.140 -0.235 6.370 1.280 ;
        RECT  2.150 -0.235 6.140 0.235 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.620 3.685 9.520 4.155 ;
        RECT  8.280 2.310 8.620 4.155 ;
        RECT  6.370 3.685 8.280 4.155 ;
        RECT  6.140 2.980 6.370 4.155 ;
        RECT  3.245 3.685 6.140 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.845 1.660 8.805 2.000 ;
        RECT  7.615 0.465 7.845 3.405 ;
        RECT  7.090 1.700 7.280 2.040 ;
        RECT  6.860 0.495 7.090 3.410 ;
        RECT  5.850 2.480 6.860 2.710 ;
        RECT  6.230 1.700 6.460 2.250 ;
        RECT  5.390 2.020 6.230 2.250 ;
        RECT  5.620 2.480 5.850 3.455 ;
        RECT  5.160 2.020 5.390 3.455 ;
        RECT  4.365 2.020 5.160 2.250 ;
        RECT  3.785 3.225 5.160 3.455 ;
        RECT  4.705 0.525 4.935 1.790 ;
        RECT  4.700 2.480 4.930 2.990 ;
        RECT  3.820 0.525 4.705 0.755 ;
        RECT  4.595 1.450 4.705 1.790 ;
        RECT  3.905 2.480 4.700 2.710 ;
        RECT  4.365 0.985 4.475 1.215 ;
        RECT  4.135 0.985 4.365 2.250 ;
        RECT  3.675 1.485 3.905 2.710 ;
        RECT  3.590 0.525 3.820 0.925 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  2.325 2.480 3.675 2.710 ;
        RECT  1.840 0.695 3.590 0.925 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 0.695 1.840 2.535 ;
        RECT  1.500 0.695 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LNCNQD1BWP7T

MACRO LNCNQD2BWP7T
    CLASS CORE ;
    FOREIGN LNCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.125 1.210 9.380 2.450 ;
        RECT  9.100 0.495 9.125 3.275 ;
        RECT  8.895 0.495 9.100 1.440 ;
        RECT  8.895 2.220 9.100 3.275 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3042 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.210 3.235 2.150 ;
        END
    END D
    PIN CDN
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.330 1.485 2.380 1.825 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 -0.235 10.080 0.235 ;
        RECT  9.615 -0.235 9.845 1.260 ;
        RECT  8.485 -0.235 9.615 0.235 ;
        RECT  8.105 -0.235 8.485 0.670 ;
        RECT  6.285 -0.235 8.105 0.235 ;
        RECT  5.935 -0.235 6.285 1.215 ;
        RECT  2.150 -0.235 5.935 0.235 ;
        RECT  1.810 -0.235 2.150 0.465 ;
        RECT  0.000 -0.235 1.810 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 3.685 10.080 4.155 ;
        RECT  9.615 2.250 9.845 4.155 ;
        RECT  8.480 3.685 9.615 4.155 ;
        RECT  8.100 3.250 8.480 4.155 ;
        RECT  6.420 3.685 8.100 4.155 ;
        RECT  6.080 3.245 6.420 4.155 ;
        RECT  3.245 3.685 6.080 4.155 ;
        RECT  3.015 3.400 3.245 4.155 ;
        RECT  1.290 3.685 3.015 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.415 1.075 8.645 3.000 ;
        RECT  7.685 1.075 8.415 1.305 ;
        RECT  7.685 2.770 8.415 3.000 ;
        RECT  7.085 1.660 7.915 2.000 ;
        RECT  7.455 0.495 7.685 1.305 ;
        RECT  7.455 2.770 7.685 3.440 ;
        RECT  6.855 0.495 7.085 3.015 ;
        RECT  6.735 0.495 6.855 1.305 ;
        RECT  5.845 2.785 6.855 3.015 ;
        RECT  6.230 1.700 6.460 2.250 ;
        RECT  5.385 2.020 6.230 2.250 ;
        RECT  5.615 2.785 5.845 3.455 ;
        RECT  5.155 2.020 5.385 3.455 ;
        RECT  4.365 2.020 5.155 2.250 ;
        RECT  3.785 3.225 5.155 3.455 ;
        RECT  4.705 0.525 4.935 1.790 ;
        RECT  4.695 2.480 4.925 2.990 ;
        RECT  3.820 0.525 4.705 0.755 ;
        RECT  4.595 1.450 4.705 1.790 ;
        RECT  3.905 2.480 4.695 2.710 ;
        RECT  4.365 0.985 4.475 1.215 ;
        RECT  4.135 0.985 4.365 2.250 ;
        RECT  3.675 1.485 3.905 2.710 ;
        RECT  3.590 0.525 3.820 0.925 ;
        RECT  3.555 2.940 3.785 3.455 ;
        RECT  2.325 2.480 3.675 2.710 ;
        RECT  1.840 0.695 3.590 0.925 ;
        RECT  2.785 2.940 3.555 3.170 ;
        RECT  2.555 2.940 2.785 3.455 ;
        RECT  2.200 3.225 2.555 3.455 ;
        RECT  2.095 2.480 2.325 2.995 ;
        RECT  0.960 2.765 2.095 2.995 ;
        RECT  1.610 0.695 1.840 2.535 ;
        RECT  1.500 0.695 1.610 1.250 ;
        RECT  1.500 2.305 1.610 2.535 ;
        RECT  0.960 1.700 1.375 2.040 ;
        RECT  0.730 0.585 0.960 2.995 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.565 0.730 2.795 ;
    END
END LNCNQD2BWP7T

MACRO LND1BWP7T
    CLASS CORE ;
    FOREIGN LND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.935 0.495 8.260 3.300 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.0040 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.580 2.415 6.700 2.645 ;
        RECT  6.580 0.485 6.645 1.305 ;
        RECT  6.415 0.485 6.580 2.645 ;
        RECT  6.300 1.115 6.415 2.645 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.405 -0.235 8.400 0.235 ;
        RECT  7.175 -0.235 7.405 1.195 ;
        RECT  5.200 -0.235 7.175 0.235 ;
        RECT  4.820 -0.235 5.200 0.670 ;
        RECT  2.420 -0.235 4.820 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.460 3.685 8.400 4.155 ;
        RECT  7.120 3.455 7.460 4.155 ;
        RECT  5.290 3.685 7.120 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.455 1.660 7.685 3.190 ;
        RECT  6.010 2.960 7.455 3.190 ;
        RECT  5.850 1.295 6.010 3.440 ;
        RECT  5.780 0.495 5.850 3.440 ;
        RECT  5.620 0.495 5.780 1.525 ;
        RECT  4.465 1.295 5.620 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.220 3.775 2.720 ;
        RECT  3.360 1.220 3.545 1.560 ;
        RECT  3.220 2.490 3.545 2.720 ;
        RECT  3.120 1.900 3.315 2.240 ;
        RECT  2.990 2.490 3.220 3.210 ;
        RECT  2.890 1.020 3.120 2.240 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  2.080 1.020 2.890 1.250 ;
        RECT  1.850 1.020 2.080 2.720 ;
        RECT  1.500 1.020 1.850 1.250 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LND1BWP7T

MACRO LND2BWP7T
    CLASS CORE ;
    FOREIGN LND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.155 9.380 2.485 ;
        RECT  8.860 1.155 9.100 1.385 ;
        RECT  8.860 2.255 9.100 2.485 ;
        RECT  8.630 0.485 8.860 1.385 ;
        RECT  8.630 2.255 8.860 3.205 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.420 1.075 7.700 2.530 ;
        RECT  7.190 0.495 7.420 1.305 ;
        RECT  7.135 2.255 7.420 2.530 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 -0.235 10.080 0.235 ;
        RECT  9.615 -0.235 9.845 1.250 ;
        RECT  8.225 -0.235 9.615 0.235 ;
        RECT  7.845 -0.235 8.225 0.820 ;
        RECT  6.715 -0.235 7.845 0.235 ;
        RECT  6.375 -0.235 6.715 1.225 ;
        RECT  5.200 -0.235 6.375 0.235 ;
        RECT  4.820 -0.235 5.200 0.670 ;
        RECT  2.420 -0.235 4.820 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 3.685 10.080 4.155 ;
        RECT  9.615 2.255 9.845 4.155 ;
        RECT  8.265 3.685 9.615 4.155 ;
        RECT  7.805 3.250 8.265 4.155 ;
        RECT  6.765 3.685 7.805 4.155 ;
        RECT  6.305 3.250 6.765 4.155 ;
        RECT  5.290 3.685 6.305 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.320 1.715 8.715 1.945 ;
        RECT  8.040 1.715 8.320 3.020 ;
        RECT  6.010 2.790 8.040 3.020 ;
        RECT  5.960 1.295 6.010 3.020 ;
        RECT  5.780 0.495 5.960 3.020 ;
        RECT  5.730 0.495 5.780 1.525 ;
        RECT  4.465 1.295 5.730 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.220 3.775 2.720 ;
        RECT  3.360 1.220 3.545 1.560 ;
        RECT  3.220 2.490 3.545 2.720 ;
        RECT  3.120 1.900 3.315 2.240 ;
        RECT  2.990 2.490 3.220 3.210 ;
        RECT  2.890 1.020 3.120 2.240 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  2.080 1.020 2.890 1.250 ;
        RECT  1.850 1.020 2.080 2.720 ;
        RECT  1.500 1.020 1.850 1.250 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LND2BWP7T

MACRO LNQD1BWP7T
    CLASS CORE ;
    FOREIGN LNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.180 7.140 2.480 ;
        RECT  6.730 1.180 6.860 1.410 ;
        RECT  6.730 2.250 6.860 2.480 ;
        RECT  6.500 0.495 6.730 1.410 ;
        RECT  6.500 2.250 6.730 3.200 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.605 -0.235 7.840 0.235 ;
        RECT  7.375 -0.235 7.605 1.235 ;
        RECT  5.360 -0.235 7.375 0.235 ;
        RECT  4.980 -0.235 5.360 0.980 ;
        RECT  2.420 -0.235 4.980 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.600 3.685 7.840 4.155 ;
        RECT  7.370 2.245 7.600 4.155 ;
        RECT  5.290 3.685 7.370 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.780 0.495 6.010 3.200 ;
        RECT  4.465 1.295 5.780 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.220 3.775 2.720 ;
        RECT  3.360 1.220 3.545 1.560 ;
        RECT  3.220 2.490 3.545 2.720 ;
        RECT  3.120 1.900 3.315 2.240 ;
        RECT  2.990 2.490 3.220 3.210 ;
        RECT  2.890 1.020 3.120 2.240 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  2.080 1.020 2.890 1.250 ;
        RECT  1.850 1.020 2.080 2.720 ;
        RECT  1.500 1.020 1.850 1.250 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LNQD1BWP7T

MACRO LNQD2BWP7T
    CLASS CORE ;
    FOREIGN LNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.445 1.180 7.700 2.480 ;
        RECT  7.420 0.495 7.445 3.200 ;
        RECT  7.215 0.495 7.420 1.410 ;
        RECT  7.215 2.250 7.420 3.200 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.3420 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.530 2.660 2.710 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.165 -0.235 8.400 0.235 ;
        RECT  7.935 -0.235 8.165 1.250 ;
        RECT  6.795 -0.235 7.935 0.235 ;
        RECT  6.415 -0.235 6.795 1.205 ;
        RECT  5.200 -0.235 6.415 0.235 ;
        RECT  4.820 -0.235 5.200 0.670 ;
        RECT  2.420 -0.235 4.820 0.235 ;
        RECT  2.080 -0.235 2.420 0.465 ;
        RECT  0.000 -0.235 2.080 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.165 3.685 8.400 4.155 ;
        RECT  7.935 2.245 8.165 4.155 ;
        RECT  6.795 3.685 7.935 4.155 ;
        RECT  6.415 2.310 6.795 4.155 ;
        RECT  5.290 3.685 6.415 4.155 ;
        RECT  5.060 2.250 5.290 4.155 ;
        RECT  2.420 3.685 5.060 4.155 ;
        RECT  2.080 3.455 2.420 4.155 ;
        RECT  1.290 3.685 2.080 4.155 ;
        RECT  0.950 3.455 1.290 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.780 0.495 6.010 3.200 ;
        RECT  4.465 1.295 5.780 1.525 ;
        RECT  4.825 1.755 5.505 1.985 ;
        RECT  4.585 1.755 4.825 3.180 ;
        RECT  4.235 1.755 4.585 1.985 ;
        RECT  3.465 2.950 4.585 3.180 ;
        RECT  3.775 2.425 4.285 2.720 ;
        RECT  4.005 0.585 4.235 1.985 ;
        RECT  3.465 0.585 4.005 0.815 ;
        RECT  3.545 1.220 3.775 2.720 ;
        RECT  3.360 1.220 3.545 1.560 ;
        RECT  3.220 2.490 3.545 2.720 ;
        RECT  3.120 1.900 3.315 2.240 ;
        RECT  2.990 2.490 3.220 3.210 ;
        RECT  2.890 1.020 3.120 2.240 ;
        RECT  0.960 2.980 2.990 3.210 ;
        RECT  2.080 1.020 2.890 1.250 ;
        RECT  1.850 1.020 2.080 2.720 ;
        RECT  1.500 1.020 1.850 1.250 ;
        RECT  1.500 2.490 1.850 2.720 ;
        RECT  0.960 1.755 1.430 1.985 ;
        RECT  0.730 0.585 0.960 3.210 ;
        RECT  0.180 0.585 0.730 0.815 ;
        RECT  0.180 2.505 0.730 2.735 ;
    END
END LNQD2BWP7T

MACRO LNSND1BWP7T
    CLASS CORE ;
    FOREIGN LNSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3033 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.615 0.495 9.940 3.185 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.075 8.820 2.535 ;
        RECT  8.405 1.075 8.540 1.305 ;
        RECT  8.120 2.305 8.540 2.535 ;
        RECT  8.175 0.485 8.405 1.305 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.2700 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 0.650 2.680 1.590 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.240 -0.235 10.080 0.235 ;
        RECT  8.780 -0.235 9.240 0.845 ;
        RECT  6.985 -0.235 8.780 0.235 ;
        RECT  6.755 -0.235 6.985 0.840 ;
        RECT  5.140 -0.235 6.755 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.250 3.685 10.080 4.155 ;
        RECT  8.790 3.250 9.250 4.155 ;
        RECT  6.800 3.685 8.790 4.155 ;
        RECT  6.455 3.445 6.800 4.155 ;
        RECT  2.545 3.685 6.455 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.135 1.660 9.365 3.020 ;
        RECT  7.035 2.790 9.135 3.020 ;
        RECT  7.710 1.590 8.310 1.935 ;
        RECT  7.430 0.500 7.710 2.560 ;
        RECT  7.290 2.330 7.430 2.560 ;
        RECT  6.805 1.160 7.035 3.020 ;
        RECT  6.480 1.160 6.805 1.390 ;
        RECT  5.980 2.790 6.805 3.020 ;
        RECT  6.250 0.605 6.480 1.390 ;
        RECT  5.990 0.605 6.250 0.835 ;
        RECT  5.750 2.790 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.935 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.675 2.705 4.875 2.935 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.375 3.225 4.295 3.455 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.275 1.070 3.760 1.300 ;
        RECT  3.165 1.685 3.530 2.050 ;
        RECT  3.135 2.940 3.375 3.455 ;
        RECT  2.060 1.820 3.165 2.050 ;
        RECT  1.455 2.940 3.135 3.170 ;
        RECT  1.830 0.935 2.060 2.710 ;
        RECT  1.760 0.935 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LNSND1BWP7T

MACRO LNSND2BWP7T
    CLASS CORE ;
    FOREIGN LNSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.2988 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.780 1.210 11.060 2.450 ;
        RECT  10.685 1.210 10.780 1.440 ;
        RECT  10.685 2.220 10.780 2.450 ;
        RECT  10.455 0.495 10.685 1.440 ;
        RECT  10.455 2.220 10.685 3.275 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.4898 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.870 0.495 9.100 1.400 ;
        RECT  8.820 2.300 9.075 2.530 ;
        RECT  8.820 1.165 8.870 1.400 ;
        RECT  8.540 1.165 8.820 2.530 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.2700 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 0.650 2.680 1.590 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.525 -0.235 11.760 0.235 ;
        RECT  11.295 -0.235 11.525 1.260 ;
        RECT  10.030 -0.235 11.295 0.235 ;
        RECT  9.650 -0.235 10.030 0.910 ;
        RECT  8.210 -0.235 9.650 0.235 ;
        RECT  7.980 -0.235 8.210 1.235 ;
        RECT  5.140 -0.235 7.980 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.520 3.685 11.760 4.155 ;
        RECT  11.290 2.250 11.520 4.155 ;
        RECT  9.925 3.685 11.290 4.155 ;
        RECT  9.545 3.250 9.925 4.155 ;
        RECT  8.355 3.685 9.545 4.155 ;
        RECT  8.015 3.250 8.355 4.155 ;
        RECT  6.880 3.685 8.015 4.155 ;
        RECT  6.485 3.455 6.880 4.155 ;
        RECT  2.545 3.685 6.485 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.975 1.620 10.205 3.020 ;
        RECT  7.060 2.790 9.975 3.020 ;
        RECT  7.710 1.655 8.290 2.030 ;
        RECT  7.430 0.585 7.710 2.530 ;
        RECT  7.075 0.585 7.430 0.815 ;
        RECT  7.290 2.300 7.430 2.530 ;
        RECT  6.830 1.110 7.060 3.020 ;
        RECT  6.670 1.110 6.830 1.340 ;
        RECT  5.980 2.790 6.830 3.020 ;
        RECT  6.440 0.605 6.670 1.340 ;
        RECT  5.990 0.605 6.440 0.835 ;
        RECT  5.750 2.790 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.935 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.655 2.705 4.875 2.935 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.405 3.225 4.295 3.455 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.245 1.070 3.760 1.300 ;
        RECT  3.165 1.685 3.530 2.050 ;
        RECT  3.165 2.940 3.405 3.455 ;
        RECT  2.060 1.820 3.165 2.050 ;
        RECT  1.455 2.940 3.165 3.170 ;
        RECT  1.830 0.730 2.060 2.710 ;
        RECT  1.760 0.730 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LNSND2BWP7T

MACRO LNSNQD1BWP7T
    CLASS CORE ;
    FOREIGN LNSNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.3033 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.5168 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.055 0.485 9.385 3.195 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.2700 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 0.650 2.680 1.590 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.520 -0.235 9.520 0.235 ;
        RECT  8.060 -0.235 8.520 1.140 ;
        RECT  6.985 -0.235 8.060 0.235 ;
        RECT  6.755 -0.235 6.985 0.840 ;
        RECT  5.140 -0.235 6.755 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.530 3.685 9.520 4.155 ;
        RECT  8.070 2.310 8.530 4.155 ;
        RECT  6.800 3.685 8.070 4.155 ;
        RECT  6.455 3.445 6.800 4.155 ;
        RECT  2.545 3.685 6.455 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.710 1.590 8.645 1.935 ;
        RECT  7.430 0.500 7.710 2.560 ;
        RECT  7.290 2.330 7.430 2.560 ;
        RECT  6.805 1.160 7.035 3.020 ;
        RECT  6.480 1.160 6.805 1.390 ;
        RECT  5.980 2.790 6.805 3.020 ;
        RECT  6.250 0.605 6.480 1.390 ;
        RECT  5.990 0.605 6.250 0.835 ;
        RECT  5.750 2.790 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.935 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.655 2.705 4.875 2.935 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.405 3.225 4.295 3.455 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.255 1.070 3.760 1.300 ;
        RECT  3.165 1.685 3.530 2.050 ;
        RECT  3.165 2.940 3.405 3.455 ;
        RECT  2.060 1.820 3.165 2.050 ;
        RECT  1.455 2.940 3.165 3.170 ;
        RECT  1.830 0.935 2.060 2.710 ;
        RECT  1.760 0.935 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LNSNQD1BWP7T

MACRO LNSNQD2BWP7T
    CLASS CORE ;
    FOREIGN LNSNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SDN
        ANTENNAGATEAREA 0.2988 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 1.700 6.170 2.150 ;
        RECT  5.740 1.210 6.020 2.150 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.4098 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.870 0.495 9.100 1.400 ;
        RECT  8.820 2.245 9.025 3.200 ;
        RECT  8.820 1.165 8.870 1.400 ;
        RECT  8.790 1.165 8.820 3.200 ;
        RECT  8.540 1.165 8.790 2.530 ;
        END
    END Q
    PIN EN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.630 1.755 0.700 2.150 ;
        END
    END EN
    PIN D
        ANTENNAGATEAREA 0.2700 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 1.210 2.825 1.590 ;
        RECT  2.380 0.650 2.680 1.590 ;
        END
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.900 -0.235 10.080 0.235 ;
        RECT  9.560 -0.235 9.900 1.180 ;
        RECT  8.210 -0.235 9.560 0.235 ;
        RECT  7.980 -0.235 8.210 1.235 ;
        RECT  5.140 -0.235 7.980 0.235 ;
        RECT  4.680 -0.235 5.140 0.885 ;
        RECT  1.285 -0.235 4.680 0.235 ;
        RECT  0.945 -0.235 1.285 0.980 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.920 3.685 10.080 4.155 ;
        RECT  9.540 2.310 9.920 4.155 ;
        RECT  8.300 3.685 9.540 4.155 ;
        RECT  8.070 2.255 8.300 4.155 ;
        RECT  6.855 3.685 8.070 4.155 ;
        RECT  6.515 2.980 6.855 4.155 ;
        RECT  2.545 3.685 6.515 4.155 ;
        RECT  2.205 3.420 2.545 4.155 ;
        RECT  1.300 3.685 2.205 4.155 ;
        RECT  0.960 3.420 1.300 4.155 ;
        RECT  0.000 3.685 0.960 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.575 1.655 8.290 2.000 ;
        RECT  7.345 0.585 7.575 3.405 ;
        RECT  7.075 0.585 7.345 0.815 ;
        RECT  6.830 1.110 7.060 2.730 ;
        RECT  6.670 1.110 6.830 1.340 ;
        RECT  5.980 2.500 6.830 2.730 ;
        RECT  6.440 0.605 6.670 1.340 ;
        RECT  5.990 0.605 6.440 0.835 ;
        RECT  5.750 2.500 5.980 3.455 ;
        RECT  4.585 3.225 5.750 3.455 ;
        RECT  5.115 1.655 5.490 1.995 ;
        RECT  4.875 1.655 5.115 2.935 ;
        RECT  4.450 1.655 4.875 1.885 ;
        RECT  3.655 2.705 4.875 2.935 ;
        RECT  4.220 0.470 4.450 1.885 ;
        RECT  3.990 2.170 4.425 2.400 ;
        RECT  3.405 3.225 4.295 3.455 ;
        RECT  3.515 0.470 4.220 0.700 ;
        RECT  3.760 1.070 3.990 2.400 ;
        RECT  3.255 1.070 3.760 1.300 ;
        RECT  3.165 1.685 3.530 2.050 ;
        RECT  3.165 2.940 3.405 3.455 ;
        RECT  2.060 1.820 3.165 2.050 ;
        RECT  1.455 2.940 3.165 3.170 ;
        RECT  1.830 0.935 2.060 2.710 ;
        RECT  1.760 0.935 1.830 1.275 ;
        RECT  1.740 2.370 1.830 2.710 ;
        RECT  1.455 1.660 1.600 2.000 ;
        RECT  1.225 1.660 1.455 3.170 ;
        RECT  0.465 2.940 1.225 3.170 ;
        RECT  0.400 0.915 0.465 1.255 ;
        RECT  0.400 2.440 0.465 3.170 ;
        RECT  0.140 0.915 0.400 3.170 ;
    END
END LNSNQD2BWP7T

MACRO MAOI222D0BWP7T
    CLASS CORE ;
    FOREIGN MAOI222D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.5229 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.950 3.780 2.905 ;
        RECT  3.210 0.950 3.500 1.190 ;
        RECT  0.935 2.675 3.500 2.905 ;
        RECT  0.695 0.925 0.935 3.310 ;
        RECT  0.180 0.925 0.695 1.155 ;
        RECT  0.180 3.080 0.695 3.310 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.365 1.260 2.710 1.540 ;
        RECT  1.770 1.260 2.365 1.765 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.915 3.000 2.375 ;
        RECT  1.540 2.135 2.770 2.375 ;
        RECT  1.220 1.210 1.540 2.375 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.895 -0.235 4.480 0.235 ;
        RECT  1.540 -0.235 1.895 0.970 ;
        RECT  0.000 -0.235 1.540 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.835 3.685 4.480 4.155 ;
        RECT  1.455 3.155 1.835 4.155 ;
        RECT  0.000 3.685 1.455 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.205 3.135 4.275 3.365 ;
        RECT  4.015 0.465 4.245 1.180 ;
        RECT  2.735 0.465 4.015 0.695 ;
        RECT  2.395 0.465 2.735 0.985 ;
    END
END MAOI222D0BWP7T

MACRO MAOI222D1BWP7T
    CLASS CORE ;
    FOREIGN MAOI222D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.4174 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.710 4.340 2.765 ;
        RECT  3.945 0.710 4.060 0.940 ;
        RECT  1.185 2.535 4.060 2.765 ;
        RECT  0.955 0.925 1.185 2.765 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.600 1.260 3.830 1.950 ;
        RECT  2.150 1.260 3.600 1.540 ;
        RECT  1.920 1.260 2.150 1.940 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.710 -0.235 4.480 0.235 ;
        RECT  2.370 -0.235 2.710 0.530 ;
        RECT  0.000 -0.235 2.370 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.785 3.685 4.480 4.155 ;
        RECT  2.435 3.455 2.785 4.155 ;
        RECT  0.000 3.685 2.435 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.895 0.775 3.585 1.005 ;
        RECT  0.465 2.995 3.580 3.225 ;
        RECT  1.565 0.465 1.895 1.005 ;
        RECT  0.180 0.465 1.565 0.695 ;
        RECT  0.235 2.405 0.465 3.225 ;
    END
END MAOI222D1BWP7T

MACRO MAOI222D2BWP7T
    CLASS CORE ;
    FOREIGN MAOI222D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.090 6.580 2.485 ;
        RECT  6.070 0.475 6.300 1.320 ;
        RECT  6.070 2.255 6.300 3.435 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 1.260 3.785 1.950 ;
        RECT  2.095 1.260 3.555 1.540 ;
        RECT  1.865 1.260 2.095 1.940 ;
        END
    END B
    PIN A
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 -0.235 7.280 0.235 ;
        RECT  6.815 -0.235 7.045 1.255 ;
        RECT  5.660 -0.235 6.815 0.235 ;
        RECT  5.280 -0.235 5.660 0.940 ;
        RECT  2.600 -0.235 5.280 0.235 ;
        RECT  2.260 -0.235 2.600 0.530 ;
        RECT  0.000 -0.235 2.260 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 3.685 7.280 4.155 ;
        RECT  6.815 2.255 7.045 4.155 ;
        RECT  5.660 3.685 6.815 4.155 ;
        RECT  5.280 2.705 5.660 4.155 ;
        RECT  2.610 3.685 5.280 4.155 ;
        RECT  2.260 3.455 2.610 4.155 ;
        RECT  0.000 3.685 2.260 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.735 1.705 6.055 1.935 ;
        RECT  5.505 1.190 5.735 2.475 ;
        RECT  4.860 1.190 5.505 1.420 ;
        RECT  4.860 2.245 5.505 2.475 ;
        RECT  4.340 1.735 5.155 1.965 ;
        RECT  4.630 0.465 4.860 1.420 ;
        RECT  4.630 2.245 4.860 3.410 ;
        RECT  4.060 0.710 4.340 2.765 ;
        RECT  3.845 0.710 4.060 0.940 ;
        RECT  1.185 2.535 4.060 2.765 ;
        RECT  1.895 0.775 3.365 1.005 ;
        RECT  0.465 2.995 3.360 3.225 ;
        RECT  1.565 0.465 1.895 1.005 ;
        RECT  0.180 0.465 1.565 0.695 ;
        RECT  0.955 0.925 1.185 2.765 ;
        RECT  0.235 2.405 0.465 3.225 ;
    END
END MAOI222D2BWP7T

MACRO MAOI22D0BWP7T
    CLASS CORE ;
    FOREIGN MAOI22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6399 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.990 3.220 2.795 ;
        RECT  2.260 0.990 2.940 1.220 ;
        RECT  2.895 2.455 2.940 2.795 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.990 1.540 1.430 1.770 ;
        RECT  0.700 1.540 0.990 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.470 1.655 3.780 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.720 2.700 2.160 ;
        RECT  2.380 1.720 2.660 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 -0.235 3.920 0.235 ;
        RECT  1.470 -0.235 1.875 0.465 ;
        RECT  0.000 -0.235 1.470 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.710 3.685 3.920 4.155 ;
        RECT  1.370 3.455 1.710 4.155 ;
        RECT  0.000 3.685 1.370 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.695 0.975 1.945 3.215 ;
        RECT  0.740 0.975 1.695 1.205 ;
        RECT  0.180 2.985 1.695 3.215 ;
    END
END MAOI22D0BWP7T

MACRO MAOI22D1BWP7T
    CLASS CORE ;
    FOREIGN MAOI22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.3717 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.110 3.780 2.740 ;
        RECT  2.770 1.110 3.500 1.340 ;
        RECT  3.240 2.510 3.500 2.740 ;
        RECT  2.425 0.465 2.770 1.340 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.675 1.540 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.030 1.610 4.340 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.675 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 -0.235 4.480 0.235 ;
        RECT  4.015 -0.235 4.245 1.245 ;
        RECT  2.030 -0.235 4.015 0.235 ;
        RECT  1.650 -0.235 2.030 0.770 ;
        RECT  0.540 -0.235 1.650 0.235 ;
        RECT  0.160 -0.235 0.540 0.930 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 3.685 4.480 4.155 ;
        RECT  1.640 2.940 2.015 4.155 ;
        RECT  0.000 3.685 1.640 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.770 3.000 4.300 3.230 ;
        RECT  2.525 2.405 2.770 3.230 ;
        RECT  1.875 1.000 2.110 2.645 ;
        RECT  1.245 1.000 1.875 1.230 ;
        RECT  0.465 2.415 1.875 2.645 ;
        RECT  0.885 0.475 1.245 1.230 ;
        RECT  0.235 2.415 0.465 3.315 ;
    END
END MAOI22D1BWP7T

MACRO MAOI22D2BWP7T
    CLASS CORE ;
    FOREIGN MAOI22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 1.170 5.460 2.665 ;
        RECT  5.180 0.495 5.205 3.435 ;
        RECT  4.975 0.495 5.180 1.400 ;
        RECT  4.975 2.375 5.180 3.435 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.615 3.780 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.505 2.805 1.845 ;
        RECT  2.380 1.505 2.660 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 -0.235 6.160 0.235 ;
        RECT  5.695 -0.235 5.925 1.245 ;
        RECT  4.580 -0.235 5.695 0.235 ;
        RECT  4.200 -0.235 4.580 1.250 ;
        RECT  1.705 -0.235 4.200 0.235 ;
        RECT  1.325 -0.235 1.705 0.865 ;
        RECT  0.000 -0.235 1.325 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 3.685 6.160 4.155 ;
        RECT  5.695 2.250 5.925 4.155 ;
        RECT  4.360 3.685 5.695 4.155 ;
        RECT  3.825 3.455 4.360 4.155 ;
        RECT  1.975 3.685 3.825 4.155 ;
        RECT  1.595 3.050 1.975 4.155 ;
        RECT  0.540 3.685 1.595 4.155 ;
        RECT  0.160 3.030 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.495 1.695 4.725 3.210 ;
        RECT  3.270 2.980 4.495 3.210 ;
        RECT  2.345 0.465 3.840 0.695 ;
        RECT  3.035 1.020 3.270 3.210 ;
        RECT  2.780 1.020 3.035 1.250 ;
        RECT  2.340 2.980 3.035 3.210 ;
        RECT  2.115 0.465 2.345 1.275 ;
        RECT  1.905 1.715 2.135 2.710 ;
        RECT  1.185 2.480 1.905 2.710 ;
        RECT  0.955 2.480 1.185 3.290 ;
        RECT  0.935 2.480 0.955 2.710 ;
        RECT  0.705 1.090 0.935 2.710 ;
        RECT  0.465 1.090 0.705 1.320 ;
        RECT  0.235 0.495 0.465 1.320 ;
    END
END MAOI22D2BWP7T

MACRO MOAI22D0BWP7T
    CLASS CORE ;
    FOREIGN MOAI22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6399 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.965 3.220 2.930 ;
        RECT  2.895 0.965 2.940 1.305 ;
        RECT  2.260 2.700 2.940 2.930 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.990 1.955 1.430 2.185 ;
        RECT  0.700 1.210 0.990 2.185 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.470 1.210 3.780 2.265 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.485 2.700 2.200 ;
        RECT  2.380 1.210 2.660 2.200 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.710 -0.235 3.920 0.235 ;
        RECT  1.370 -0.235 1.710 0.465 ;
        RECT  0.000 -0.235 1.370 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 3.685 3.920 4.155 ;
        RECT  1.470 3.455 1.875 4.155 ;
        RECT  0.000 3.685 1.470 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.695 0.705 1.945 2.945 ;
        RECT  0.180 0.705 1.695 0.935 ;
        RECT  0.740 2.715 1.695 2.945 ;
    END
END MOAI22D0BWP7T

MACRO MOAI22D1BWP7T
    CLASS CORE ;
    FOREIGN MOAI22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.095 3.780 3.280 ;
        RECT  3.365 1.095 3.500 1.325 ;
        RECT  2.545 3.050 3.500 3.280 ;
        RECT  3.025 1.020 3.365 1.325 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.655 1.540 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.670 0.800 1.900 ;
        RECT  0.140 1.670 0.420 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.030 1.210 4.340 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.610 3.220 2.750 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.930 -0.235 4.480 0.235 ;
        RECT  1.550 -0.235 1.930 0.805 ;
        RECT  0.000 -0.235 1.550 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.240 3.685 4.480 4.155 ;
        RECT  4.010 2.520 4.240 4.155 ;
        RECT  2.175 3.685 4.010 4.155 ;
        RECT  1.735 3.455 2.175 4.155 ;
        RECT  0.640 3.685 1.735 4.155 ;
        RECT  0.260 3.115 0.640 4.155 ;
        RECT  0.000 3.685 0.260 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.800 0.465 4.030 0.860 ;
        RECT  2.590 0.465 3.800 0.695 ;
        RECT  2.360 0.465 2.590 1.305 ;
        RECT  2.125 1.670 2.290 2.010 ;
        RECT  2.115 1.110 2.125 2.010 ;
        RECT  1.885 1.110 2.115 3.225 ;
        RECT  0.550 1.110 1.885 1.340 ;
        RECT  0.985 2.995 1.885 3.225 ;
        RECT  0.320 0.495 0.550 1.340 ;
    END
END MOAI22D1BWP7T

MACRO MOAI22D2BWP7T
    CLASS CORE ;
    FOREIGN MOAI22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.3398 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.200 1.170 5.460 2.710 ;
        RECT  5.180 1.170 5.200 3.400 ;
        RECT  5.160 1.170 5.180 1.400 ;
        RECT  4.970 2.375 5.180 3.400 ;
        RECT  4.930 0.495 5.160 1.400 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.825 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.365 1.575 3.220 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.640 1.405 2.150 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.920 -0.235 6.160 0.235 ;
        RECT  5.690 -0.235 5.920 1.260 ;
        RECT  4.315 -0.235 5.690 0.235 ;
        RECT  3.945 -0.235 4.315 0.465 ;
        RECT  2.015 -0.235 3.945 0.235 ;
        RECT  1.655 -0.235 2.015 0.465 ;
        RECT  0.545 -0.235 1.655 0.235 ;
        RECT  0.165 -0.235 0.545 0.960 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.920 3.685 6.160 4.155 ;
        RECT  5.690 2.255 5.920 4.155 ;
        RECT  4.475 3.685 5.690 4.155 ;
        RECT  4.110 3.455 4.475 4.155 ;
        RECT  1.675 3.685 4.110 4.155 ;
        RECT  1.425 2.975 1.675 4.155 ;
        RECT  0.000 3.685 1.425 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.515 1.655 4.795 1.885 ;
        RECT  4.500 0.715 4.515 1.885 ;
        RECT  4.270 0.715 4.500 3.205 ;
        RECT  2.425 0.715 4.270 0.945 ;
        RECT  2.845 2.975 4.270 3.205 ;
        RECT  2.425 2.445 3.925 2.675 ;
        RECT  2.195 2.445 2.425 3.390 ;
        RECT  1.900 1.640 2.095 1.980 ;
        RECT  1.670 0.710 1.900 2.680 ;
        RECT  0.900 0.710 1.670 0.940 ;
        RECT  1.065 2.450 1.670 2.680 ;
        RECT  0.825 2.450 1.065 3.170 ;
        RECT  0.465 2.940 0.825 3.170 ;
        RECT  0.235 2.940 0.465 3.440 ;
    END
END MOAI22D2BWP7T

MACRO MUX2D0BWP7T
    CLASS CORE ;
    FOREIGN MUX2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.570 0.570 4.900 3.095 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 1.150 2.805 1.490 ;
        RECT  0.980 1.150 2.575 1.380 ;
        RECT  0.700 1.150 0.980 2.150 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 3.785 2.710 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.750 2.100 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 -0.235 5.040 0.235 ;
        RECT  3.760 -0.235 4.100 0.785 ;
        RECT  1.285 -0.235 3.760 0.235 ;
        RECT  0.905 -0.235 1.285 0.805 ;
        RECT  0.000 -0.235 0.905 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 3.685 5.040 4.155 ;
        RECT  3.760 2.940 4.100 4.155 ;
        RECT  1.260 3.685 3.760 4.155 ;
        RECT  0.920 2.840 1.260 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.095 1.020 4.325 1.560 ;
        RECT  3.270 1.020 4.095 1.280 ;
        RECT  3.040 0.600 3.270 3.090 ;
        RECT  2.300 0.600 3.040 0.830 ;
        RECT  2.340 2.860 3.040 3.090 ;
        RECT  2.520 1.865 2.750 2.610 ;
        RECT  0.480 2.380 2.520 2.610 ;
        RECT  0.470 2.380 0.480 2.975 ;
        RECT  0.240 0.570 0.470 2.975 ;
    END
END MUX2D0BWP7T

MACRO MUX2D1BWP7T
    CLASS CORE ;
    FOREIGN MUX2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.810 1.210 4.900 2.150 ;
        RECT  4.570 0.465 4.810 3.270 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.150 2.750 1.540 ;
        RECT  0.980 1.260 2.520 1.540 ;
        RECT  0.700 1.260 0.980 2.150 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 1.660 3.780 2.710 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.100 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 -0.235 5.040 0.235 ;
        RECT  3.760 -0.235 4.100 0.670 ;
        RECT  1.260 -0.235 3.760 0.235 ;
        RECT  0.920 -0.235 1.260 0.680 ;
        RECT  0.000 -0.235 0.920 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.125 3.685 5.040 4.155 ;
        RECT  3.745 2.940 4.125 4.155 ;
        RECT  1.260 3.685 3.745 4.155 ;
        RECT  0.920 2.940 1.260 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.110 0.900 4.340 1.945 ;
        RECT  3.215 0.900 4.110 1.160 ;
        RECT  3.210 0.490 3.215 1.160 ;
        RECT  2.980 0.490 3.210 3.080 ;
        RECT  2.300 0.490 2.980 0.720 ;
        RECT  2.340 2.850 2.980 3.080 ;
        RECT  2.520 1.850 2.750 2.610 ;
        RECT  2.055 2.380 2.520 2.610 ;
        RECT  1.805 2.380 2.055 2.710 ;
        RECT  0.480 2.480 1.805 2.710 ;
        RECT  0.470 2.480 0.480 3.085 ;
        RECT  0.240 0.465 0.470 3.085 ;
    END
END MUX2D1BWP7T

MACRO MUX2D2BWP7T
    CLASS CORE ;
    FOREIGN MUX2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.710 0.780 4.900 2.710 ;
        RECT  4.620 0.780 4.710 3.255 ;
        RECT  4.360 0.780 4.620 1.020 ;
        RECT  4.410 2.445 4.620 3.255 ;
        END
    END Z
    PIN S
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.150 2.750 1.540 ;
        RECT  0.980 1.260 2.520 1.540 ;
        RECT  0.700 1.260 0.980 2.150 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.470 1.725 3.780 2.710 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.100 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.370 -0.235 5.600 0.235 ;
        RECT  5.130 -0.235 5.370 1.250 ;
        RECT  3.980 -0.235 5.130 0.235 ;
        RECT  3.640 -0.235 3.980 0.950 ;
        RECT  1.260 -0.235 3.640 0.235 ;
        RECT  0.920 -0.235 1.260 0.680 ;
        RECT  0.000 -0.235 0.920 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.370 3.685 5.600 4.155 ;
        RECT  5.130 2.255 5.370 4.155 ;
        RECT  4.005 3.685 5.130 4.155 ;
        RECT  3.625 2.940 4.005 4.155 ;
        RECT  1.295 3.685 3.625 4.155 ;
        RECT  0.915 2.940 1.295 4.155 ;
        RECT  0.000 3.685 0.915 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.160 1.260 4.390 1.945 ;
        RECT  3.245 1.260 4.160 1.490 ;
        RECT  3.240 0.490 3.245 1.490 ;
        RECT  2.980 0.490 3.240 3.180 ;
        RECT  2.300 0.490 2.980 0.720 ;
        RECT  2.320 2.950 2.980 3.180 ;
        RECT  2.500 1.850 2.740 2.710 ;
        RECT  0.480 2.480 2.500 2.710 ;
        RECT  0.470 2.480 0.480 3.085 ;
        RECT  0.240 0.465 0.470 3.085 ;
    END
END MUX2D2BWP7T

MACRO MUX2ND0BWP7T
    CLASS CORE ;
    FOREIGN MUX2ND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6947 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.150 4.340 3.000 ;
        RECT  3.505 1.150 4.060 1.380 ;
        RECT  3.455 2.770 4.060 3.000 ;
        RECT  3.275 0.495 3.505 1.380 ;
        RECT  3.225 2.770 3.455 3.110 ;
        RECT  2.285 0.495 3.275 0.725 ;
        RECT  2.325 2.880 3.225 3.110 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.125 2.865 1.355 ;
        RECT  0.700 1.125 0.980 2.150 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 3.780 2.150 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.755 2.100 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.170 -0.235 4.480 0.235 ;
        RECT  3.790 -0.235 4.170 0.875 ;
        RECT  1.315 -0.235 3.790 0.235 ;
        RECT  0.850 -0.235 1.315 0.710 ;
        RECT  0.000 -0.235 0.850 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.180 3.685 4.480 4.155 ;
        RECT  3.800 3.250 4.180 4.155 ;
        RECT  1.265 3.685 3.800 4.155 ;
        RECT  0.885 2.995 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.470 1.770 2.710 2.610 ;
        RECT  1.940 2.380 2.470 2.610 ;
        RECT  1.710 2.380 1.940 2.680 ;
        RECT  0.465 2.450 1.710 2.680 ;
        RECT  0.235 0.465 0.465 3.200 ;
    END
END MUX2ND0BWP7T

MACRO MUX2ND1BWP7T
    CLASS CORE ;
    FOREIGN MUX2ND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.695 0.490 6.020 3.290 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 1.070 2.735 1.410 ;
        RECT  0.980 1.070 2.475 1.300 ;
        RECT  0.700 1.070 0.980 2.150 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 1.260 3.830 2.100 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.600 2.100 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.220 -0.235 6.160 0.235 ;
        RECT  4.880 -0.235 5.220 0.470 ;
        RECT  3.955 -0.235 4.880 0.235 ;
        RECT  3.575 -0.235 3.955 0.715 ;
        RECT  1.270 -0.235 3.575 0.235 ;
        RECT  0.890 -0.235 1.270 0.710 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.255 3.685 6.160 4.155 ;
        RECT  4.875 3.455 5.255 4.155 ;
        RECT  3.955 3.685 4.875 4.155 ;
        RECT  3.575 2.940 3.955 4.155 ;
        RECT  1.265 3.685 3.575 4.155 ;
        RECT  0.885 2.920 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.990 0.930 5.220 3.025 ;
        RECT  4.380 0.930 4.990 1.170 ;
        RECT  4.310 2.795 4.990 3.025 ;
        RECT  4.305 1.935 4.430 2.165 ;
        RECT  4.075 1.935 4.305 2.565 ;
        RECT  3.210 2.335 4.075 2.565 ;
        RECT  2.980 0.495 3.210 3.160 ;
        RECT  2.260 0.495 2.980 0.725 ;
        RECT  2.270 2.930 2.980 3.160 ;
        RECT  2.435 1.740 2.675 2.680 ;
        RECT  0.465 2.450 2.435 2.680 ;
        RECT  0.235 0.465 0.465 3.090 ;
    END
END MUX2ND1BWP7T

MACRO MUX2ND2BWP7T
    CLASS CORE ;
    FOREIGN MUX2ND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.325 1.060 6.580 2.710 ;
        RECT  6.300 0.475 6.325 3.265 ;
        RECT  6.095 0.475 6.300 1.290 ;
        RECT  6.095 2.435 6.300 3.265 ;
        END
    END ZN
    PIN S
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.070 2.790 1.540 ;
        RECT  0.945 1.260 2.560 1.540 ;
        RECT  0.715 1.260 0.945 2.000 ;
        END
    END S
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.680 3.855 2.710 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3492 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 1.820 2.150 2.100 ;
        RECT  1.350 1.780 1.690 2.100 ;
        RECT  1.210 1.820 1.350 2.100 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.050 -0.235 7.280 0.235 ;
        RECT  6.810 -0.235 7.050 1.270 ;
        RECT  5.660 -0.235 6.810 0.235 ;
        RECT  5.320 -0.235 5.660 0.970 ;
        RECT  4.100 -0.235 5.320 0.235 ;
        RECT  3.760 -0.235 4.100 0.845 ;
        RECT  1.280 -0.235 3.760 0.235 ;
        RECT  0.900 -0.235 1.280 0.710 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.050 3.685 7.280 4.155 ;
        RECT  6.810 2.255 7.050 4.155 ;
        RECT  5.660 3.685 6.810 4.155 ;
        RECT  5.320 2.775 5.660 4.155 ;
        RECT  4.125 3.685 5.320 4.155 ;
        RECT  3.745 3.065 4.125 4.155 ;
        RECT  1.265 3.685 3.745 4.155 ;
        RECT  0.925 2.820 1.265 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.390 1.320 5.620 2.515 ;
        RECT  4.805 1.320 5.390 1.550 ;
        RECT  4.770 2.285 5.390 2.515 ;
        RECT  4.575 0.650 4.805 1.550 ;
        RECT  4.530 2.285 4.770 3.310 ;
        RECT  4.315 1.780 4.600 2.010 ;
        RECT  4.085 1.150 4.315 2.010 ;
        RECT  3.250 1.150 4.085 1.380 ;
        RECT  3.020 0.495 3.250 3.050 ;
        RECT  2.315 0.495 3.020 0.725 ;
        RECT  2.360 2.820 3.020 3.050 ;
        RECT  2.545 1.770 2.785 2.580 ;
        RECT  0.465 2.350 2.545 2.580 ;
        RECT  0.235 0.465 0.465 2.960 ;
    END
END MUX2ND2BWP7T

MACRO MUX3D0BWP7T
    CLASS CORE ;
    FOREIGN MUX3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.165 1.210 8.260 2.150 ;
        RECT  7.935 0.945 8.165 3.130 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.390 1.550 4.435 1.890 ;
        RECT  4.010 1.260 4.390 2.100 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 2.465 2.400 2.695 ;
        RECT  1.770 2.465 2.000 3.205 ;
        RECT  0.980 2.975 1.770 3.205 ;
        RECT  0.750 1.770 0.980 3.205 ;
        RECT  0.615 1.770 0.750 2.710 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.785 1.650 7.140 2.710 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.485 -0.235 8.400 0.235 ;
        RECT  7.105 -0.235 7.485 0.940 ;
        RECT  3.960 -0.235 7.105 0.235 ;
        RECT  3.620 -0.235 3.960 0.845 ;
        RECT  1.265 -0.235 3.620 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.530 3.685 8.400 4.155 ;
        RECT  7.145 2.940 7.530 4.155 ;
        RECT  3.975 3.685 7.145 4.155 ;
        RECT  3.595 3.250 3.975 4.155 ;
        RECT  1.305 3.685 3.595 4.155 ;
        RECT  0.925 3.455 1.305 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.455 1.170 7.685 1.985 ;
        RECT  6.105 1.170 7.455 1.400 ;
        RECT  5.875 0.965 6.105 3.055 ;
        RECT  5.405 0.995 5.635 3.020 ;
        RECT  5.385 0.995 5.405 1.225 ;
        RECT  3.100 2.790 5.405 3.020 ;
        RECT  5.155 0.885 5.385 1.225 ;
        RECT  4.895 1.770 5.160 2.000 ;
        RECT  4.665 0.665 4.895 2.560 ;
        RECT  4.390 0.665 4.665 0.895 ;
        RECT  4.390 2.330 4.665 2.560 ;
        RECT  2.870 0.650 3.100 3.440 ;
        RECT  2.300 0.650 2.870 0.880 ;
        RECT  2.300 3.210 2.870 3.440 ;
        RECT  2.085 1.130 2.315 1.970 ;
        RECT  0.465 1.130 2.085 1.360 ;
        RECT  0.380 3.110 0.520 3.340 ;
        RECT  0.380 0.575 0.465 1.360 ;
        RECT  0.235 0.575 0.380 3.340 ;
        RECT  0.150 1.130 0.235 3.340 ;
    END
END MUX3D0BWP7T

MACRO MUX3D1BWP7T
    CLASS CORE ;
    FOREIGN MUX3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.165 1.210 8.260 2.150 ;
        RECT  7.935 0.475 8.165 3.385 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.390 1.550 4.435 1.890 ;
        RECT  4.010 1.260 4.390 2.100 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 2.465 2.400 2.695 ;
        RECT  1.770 2.465 2.000 3.205 ;
        RECT  0.980 2.975 1.770 3.205 ;
        RECT  0.750 1.770 0.980 3.205 ;
        RECT  0.615 1.770 0.750 2.710 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.785 1.650 7.140 2.710 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3483 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.525 -0.235 8.400 0.235 ;
        RECT  7.145 -0.235 7.525 0.930 ;
        RECT  3.960 -0.235 7.145 0.235 ;
        RECT  3.620 -0.235 3.960 0.670 ;
        RECT  1.265 -0.235 3.620 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.530 3.685 8.400 4.155 ;
        RECT  7.145 2.940 7.530 4.155 ;
        RECT  3.975 3.685 7.145 4.155 ;
        RECT  3.595 3.250 3.975 4.155 ;
        RECT  1.305 3.685 3.595 4.155 ;
        RECT  0.925 3.455 1.305 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.455 1.170 7.685 1.985 ;
        RECT  6.105 1.170 7.455 1.400 ;
        RECT  5.875 0.965 6.105 3.310 ;
        RECT  5.405 0.995 5.635 3.020 ;
        RECT  5.385 0.995 5.405 1.225 ;
        RECT  5.385 2.790 5.405 3.020 ;
        RECT  5.155 0.885 5.385 1.225 ;
        RECT  5.155 2.790 5.385 3.330 ;
        RECT  4.895 1.780 5.160 2.010 ;
        RECT  3.100 2.790 5.155 3.020 ;
        RECT  4.665 0.585 4.895 2.560 ;
        RECT  4.390 0.585 4.665 0.815 ;
        RECT  4.390 2.330 4.665 2.560 ;
        RECT  2.870 0.550 3.100 3.440 ;
        RECT  2.300 0.550 2.870 0.780 ;
        RECT  2.300 3.210 2.870 3.440 ;
        RECT  2.085 1.055 2.315 1.970 ;
        RECT  0.465 1.055 2.085 1.285 ;
        RECT  0.380 3.110 0.520 3.340 ;
        RECT  0.380 0.575 0.465 1.285 ;
        RECT  0.235 0.575 0.380 3.340 ;
        RECT  0.150 1.055 0.235 3.340 ;
    END
END MUX3D1BWP7T

MACRO MUX3D2BWP7T
    CLASS CORE ;
    FOREIGN MUX3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.005 0.650 8.260 2.710 ;
        RECT  7.980 0.475 8.005 3.385 ;
        RECT  7.775 0.475 7.980 0.880 ;
        RECT  7.775 2.310 7.980 3.385 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.5688 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 1.140 4.340 2.150 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.4635 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.650 1.105 2.810 1.445 ;
        RECT  2.420 1.105 2.650 2.610 ;
        RECT  2.000 2.380 2.420 2.610 ;
        RECT  1.770 2.380 2.000 3.205 ;
        RECT  0.980 2.975 1.770 3.205 ;
        RECT  0.750 1.760 0.980 3.205 ;
        RECT  0.600 1.760 0.750 2.710 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.4131 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.815 1.725 7.140 2.710 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.670 1.540 2.710 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.725 -0.235 8.960 0.235 ;
        RECT  8.495 -0.235 8.725 1.225 ;
        RECT  7.365 -0.235 8.495 0.235 ;
        RECT  6.985 -0.235 7.365 0.930 ;
        RECT  3.960 -0.235 6.985 0.235 ;
        RECT  3.620 -0.235 3.960 0.670 ;
        RECT  1.265 -0.235 3.620 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.725 3.685 8.960 4.155 ;
        RECT  8.495 2.255 8.725 4.155 ;
        RECT  7.370 3.685 8.495 4.155 ;
        RECT  6.985 2.940 7.370 4.155 ;
        RECT  4.000 3.685 6.985 4.155 ;
        RECT  3.660 3.455 4.000 4.155 ;
        RECT  1.305 3.685 3.660 4.155 ;
        RECT  0.925 3.455 1.305 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.500 1.170 7.730 1.985 ;
        RECT  6.105 1.170 7.500 1.400 ;
        RECT  5.875 0.965 6.105 3.310 ;
        RECT  5.415 0.995 5.645 3.225 ;
        RECT  5.385 0.995 5.415 1.225 ;
        RECT  3.270 2.995 5.415 3.225 ;
        RECT  5.155 0.885 5.385 1.225 ;
        RECT  4.860 1.780 5.185 2.120 ;
        RECT  4.630 0.585 4.860 2.610 ;
        RECT  4.390 0.585 4.630 0.815 ;
        RECT  4.390 2.380 4.630 2.610 ;
        RECT  3.040 0.550 3.270 3.440 ;
        RECT  2.300 0.550 3.040 0.780 ;
        RECT  2.300 3.210 3.040 3.440 ;
        RECT  1.945 1.055 2.175 1.995 ;
        RECT  0.465 1.055 1.945 1.285 ;
        RECT  0.365 3.110 0.520 3.340 ;
        RECT  0.365 0.575 0.465 1.285 ;
        RECT  0.235 0.575 0.365 3.340 ;
        RECT  0.135 1.055 0.235 3.340 ;
    END
END MUX3D2BWP7T

MACRO MUX3ND0BWP7T
    CLASS CORE ;
    FOREIGN MUX3ND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.840 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.7702 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.210 6.580 2.710 ;
        RECT  6.175 1.210 6.300 1.440 ;
        RECT  6.175 2.480 6.300 2.710 ;
        RECT  5.945 0.965 6.175 1.440 ;
        RECT  5.945 2.480 6.175 3.055 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.390 1.550 4.435 1.890 ;
        RECT  4.010 1.260 4.390 2.100 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 2.465 2.400 2.695 ;
        RECT  1.770 2.465 2.000 3.205 ;
        RECT  0.980 2.975 1.770 3.205 ;
        RECT  0.750 1.770 0.980 3.205 ;
        RECT  0.615 1.770 0.750 2.710 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.650 7.140 2.710 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2430 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.605 -0.235 7.840 0.235 ;
        RECT  7.375 -0.235 7.605 1.265 ;
        RECT  3.960 -0.235 7.375 0.235 ;
        RECT  3.620 -0.235 3.960 0.765 ;
        RECT  1.265 -0.235 3.620 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.605 3.685 7.840 4.155 ;
        RECT  7.375 2.725 7.605 4.155 ;
        RECT  3.975 3.685 7.375 4.155 ;
        RECT  3.595 3.250 3.975 4.155 ;
        RECT  1.305 3.685 3.595 4.155 ;
        RECT  0.925 3.455 1.305 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.405 0.995 5.635 3.020 ;
        RECT  5.385 0.995 5.405 1.225 ;
        RECT  3.100 2.790 5.405 3.020 ;
        RECT  5.155 0.885 5.385 1.225 ;
        RECT  4.895 1.770 5.160 2.000 ;
        RECT  4.665 0.585 4.895 2.560 ;
        RECT  4.390 0.585 4.665 0.815 ;
        RECT  4.390 2.330 4.665 2.560 ;
        RECT  2.870 0.570 3.100 3.440 ;
        RECT  2.300 0.570 2.870 0.800 ;
        RECT  2.300 3.210 2.870 3.440 ;
        RECT  2.085 1.055 2.315 1.970 ;
        RECT  0.465 1.055 2.085 1.285 ;
        RECT  0.380 3.110 0.520 3.340 ;
        RECT  0.380 0.575 0.465 1.285 ;
        RECT  0.235 0.575 0.380 3.340 ;
        RECT  0.150 1.055 0.235 3.340 ;
    END
END MUX3ND0BWP7T

MACRO MUX3ND1BWP7T
    CLASS CORE ;
    FOREIGN MUX3ND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.285 1.035 9.380 2.470 ;
        RECT  9.100 0.465 9.285 3.285 ;
        RECT  9.055 0.465 9.100 1.275 ;
        RECT  9.055 2.250 9.100 3.285 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.890 1.145 4.120 1.540 ;
        RECT  2.890 1.260 3.890 1.540 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 2.410 2.345 2.750 ;
        RECT  1.770 2.410 2.000 3.205 ;
        RECT  0.980 2.975 1.770 3.205 ;
        RECT  0.750 1.770 0.980 3.205 ;
        RECT  0.580 1.770 0.750 2.710 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.580 1.705 6.945 1.935 ;
        RECT  6.300 1.705 6.580 2.710 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 3.780 2.710 ;
        RECT  3.160 1.770 3.500 2.010 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3483 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.565 -0.235 9.520 0.235 ;
        RECT  8.335 -0.235 8.565 0.725 ;
        RECT  7.275 -0.235 8.335 0.235 ;
        RECT  6.895 -0.235 7.275 0.930 ;
        RECT  3.815 -0.235 6.895 0.235 ;
        RECT  3.475 -0.235 3.815 0.825 ;
        RECT  1.265 -0.235 3.475 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.565 3.685 9.520 4.155 ;
        RECT  8.335 3.090 8.565 4.155 ;
        RECT  7.390 3.685 8.335 4.155 ;
        RECT  7.005 2.940 7.390 4.155 ;
        RECT  4.010 3.685 7.005 4.155 ;
        RECT  3.670 3.455 4.010 4.155 ;
        RECT  1.305 3.685 3.670 4.155 ;
        RECT  0.925 3.455 1.305 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.025 1.715 8.760 1.945 ;
        RECT  8.020 1.715 8.025 2.650 ;
        RECT  7.790 0.965 8.020 2.650 ;
        RECT  7.685 0.965 7.790 1.305 ;
        RECT  7.405 1.645 7.560 1.985 ;
        RECT  7.175 1.170 7.405 1.985 ;
        RECT  5.875 1.170 7.175 1.400 ;
        RECT  5.875 3.025 6.035 3.255 ;
        RECT  5.645 0.965 5.875 3.255 ;
        RECT  5.260 1.120 5.405 3.210 ;
        RECT  5.175 1.120 5.260 3.455 ;
        RECT  5.155 1.120 5.175 1.350 ;
        RECT  5.030 2.980 5.175 3.455 ;
        RECT  4.925 1.010 5.155 1.350 ;
        RECT  2.805 2.980 5.030 3.210 ;
        RECT  4.730 1.715 4.920 2.055 ;
        RECT  4.695 1.715 4.730 2.605 ;
        RECT  4.465 0.515 4.695 2.605 ;
        RECT  4.195 0.515 4.465 0.745 ;
        RECT  4.390 2.375 4.465 2.605 ;
        RECT  2.660 1.955 2.805 3.440 ;
        RECT  2.575 0.550 2.660 3.440 ;
        RECT  2.430 0.550 2.575 2.185 ;
        RECT  2.300 3.210 2.575 3.440 ;
        RECT  2.155 0.550 2.430 0.780 ;
        RECT  1.970 1.055 2.200 1.920 ;
        RECT  0.465 1.055 1.970 1.285 ;
        RECT  0.350 3.110 0.520 3.340 ;
        RECT  0.350 0.575 0.465 1.285 ;
        RECT  0.235 0.575 0.350 3.340 ;
        RECT  0.120 1.055 0.235 3.340 ;
    END
END MUX3ND1BWP7T

MACRO MUX3ND2BWP7T
    CLASS CORE ;
    FOREIGN MUX3ND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.685 1.210 9.940 2.710 ;
        RECT  9.660 0.465 9.685 3.285 ;
        RECT  9.455 0.465 9.660 1.450 ;
        RECT  9.455 2.460 9.660 3.285 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.5535 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.890 1.145 4.120 1.540 ;
        RECT  2.890 1.260 3.890 1.540 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.5247 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 2.255 2.345 2.595 ;
        RECT  1.770 2.255 2.000 3.205 ;
        RECT  0.980 2.975 1.770 3.205 ;
        RECT  0.750 1.770 0.980 3.205 ;
        RECT  0.580 1.770 0.750 2.710 ;
        END
    END S0
    PIN I2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.650 7.140 2.710 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 3.780 2.710 ;
        RECT  3.160 1.770 3.500 2.010 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.3483 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 -0.235 10.640 0.235 ;
        RECT  10.175 -0.235 10.405 1.195 ;
        RECT  8.965 -0.235 10.175 0.235 ;
        RECT  8.735 -0.235 8.965 1.195 ;
        RECT  7.625 -0.235 8.735 0.235 ;
        RECT  7.245 -0.235 7.625 0.930 ;
        RECT  3.815 -0.235 7.245 0.235 ;
        RECT  3.475 -0.235 3.815 0.825 ;
        RECT  1.265 -0.235 3.475 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 3.685 10.640 4.155 ;
        RECT  10.175 2.255 10.405 4.155 ;
        RECT  8.965 3.685 10.175 4.155 ;
        RECT  8.735 2.255 8.965 4.155 ;
        RECT  7.545 3.685 8.735 4.155 ;
        RECT  7.315 2.920 7.545 4.155 ;
        RECT  4.010 3.685 7.315 4.155 ;
        RECT  3.670 3.400 4.010 4.155 ;
        RECT  1.305 3.685 3.670 4.155 ;
        RECT  0.925 3.455 1.305 4.155 ;
        RECT  0.000 3.685 0.925 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.265 1.715 9.160 1.945 ;
        RECT  8.030 0.495 8.265 3.315 ;
        RECT  7.645 1.645 7.800 1.985 ;
        RECT  7.415 1.170 7.645 1.985 ;
        RECT  6.115 1.170 7.415 1.400 ;
        RECT  6.115 3.025 6.275 3.255 ;
        RECT  5.885 0.965 6.115 3.255 ;
        RECT  5.415 1.120 5.645 3.170 ;
        RECT  5.395 1.120 5.415 1.350 ;
        RECT  2.805 2.940 5.415 3.170 ;
        RECT  5.165 1.010 5.395 1.350 ;
        RECT  4.795 1.715 4.985 2.055 ;
        RECT  4.760 1.715 4.795 2.645 ;
        RECT  4.530 0.515 4.760 2.645 ;
        RECT  4.260 0.515 4.530 0.745 ;
        RECT  4.455 2.415 4.530 2.645 ;
        RECT  2.660 1.780 2.805 3.440 ;
        RECT  2.575 0.550 2.660 3.440 ;
        RECT  2.430 0.550 2.575 2.010 ;
        RECT  2.300 3.210 2.575 3.440 ;
        RECT  2.155 0.550 2.430 0.780 ;
        RECT  1.970 1.055 2.200 1.920 ;
        RECT  0.465 1.055 1.970 1.285 ;
        RECT  0.350 3.110 0.520 3.340 ;
        RECT  0.350 0.575 0.465 1.285 ;
        RECT  0.235 0.575 0.350 3.340 ;
        RECT  0.120 1.055 0.235 3.340 ;
    END
END MUX3ND2BWP7T

MACRO MUX4D0BWP7T
    CLASS CORE ;
    FOREIGN MUX4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.735 0.940 11.060 2.925 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 1.260 6.890 2.065 ;
        RECT  5.690 1.260 6.660 1.540 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.6399 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.170 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 2.020 6.265 2.250 ;
        RECT  5.740 1.770 6.020 2.710 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.365 1.820 4.950 2.100 ;
        RECT  4.010 1.780 4.365 2.100 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        RECT  1.245 1.770 1.260 2.140 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 1.770 3.780 2.150 ;
        RECT  3.355 1.770 3.695 2.265 ;
        RECT  2.940 1.770 3.355 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.295 -0.235 11.200 0.235 ;
        RECT  9.955 -0.235 10.295 1.150 ;
        RECT  6.665 -0.235 9.955 0.235 ;
        RECT  6.325 -0.235 6.665 0.465 ;
        RECT  4.105 -0.235 6.325 0.235 ;
        RECT  3.765 -0.235 4.105 0.740 ;
        RECT  1.240 -0.235 3.765 0.235 ;
        RECT  0.900 -0.235 1.240 1.080 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 3.685 11.200 4.155 ;
        RECT  9.960 2.770 10.300 4.155 ;
        RECT  6.465 3.685 9.960 4.155 ;
        RECT  6.125 3.455 6.465 4.155 ;
        RECT  3.975 3.685 6.125 4.155 ;
        RECT  3.635 3.050 3.975 4.155 ;
        RECT  1.240 3.685 3.635 4.155 ;
        RECT  0.900 3.250 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.235 1.380 10.465 2.540 ;
        RECT  9.540 1.380 10.235 1.610 ;
        RECT  9.545 2.310 10.235 2.540 ;
        RECT  8.810 1.850 10.005 2.080 ;
        RECT  9.315 2.310 9.545 3.345 ;
        RECT  9.310 0.870 9.540 1.610 ;
        RECT  6.915 3.115 9.315 3.345 ;
        RECT  8.580 0.900 8.810 2.825 ;
        RECT  7.860 0.705 8.090 2.825 ;
        RECT  5.460 0.705 7.860 0.935 ;
        RECT  7.400 1.275 7.630 2.715 ;
        RECT  7.370 1.275 7.400 1.505 ;
        RECT  7.370 2.485 7.400 2.715 ;
        RECT  7.140 1.165 7.370 1.505 ;
        RECT  7.140 2.485 7.370 2.825 ;
        RECT  6.685 2.940 6.915 3.345 ;
        RECT  5.635 2.940 6.685 3.170 ;
        RECT  5.405 2.940 5.635 3.285 ;
        RECT  5.230 0.705 5.460 2.675 ;
        RECT  4.710 3.055 5.405 3.285 ;
        RECT  5.035 1.220 5.230 1.450 ;
        RECT  5.190 2.420 5.230 2.675 ;
        RECT  4.960 2.420 5.190 2.825 ;
        RECT  4.770 0.605 5.000 0.945 ;
        RECT  4.570 0.715 4.770 0.945 ;
        RECT  4.475 2.590 4.710 3.285 ;
        RECT  4.340 0.715 4.570 1.200 ;
        RECT  2.635 2.590 4.475 2.820 ;
        RECT  3.145 0.970 4.340 1.200 ;
        RECT  2.905 0.660 3.145 1.200 ;
        RECT  2.000 0.660 2.905 0.890 ;
        RECT  2.405 1.165 2.635 3.225 ;
        RECT  2.230 2.885 2.405 3.225 ;
        RECT  2.000 2.205 2.145 2.545 ;
        RECT  1.770 0.660 2.000 2.545 ;
        RECT  0.465 1.310 1.770 1.540 ;
        RECT  0.345 3.110 0.520 3.340 ;
        RECT  0.345 0.840 0.465 1.540 ;
        RECT  0.235 0.840 0.345 3.340 ;
        RECT  0.115 1.310 0.235 3.340 ;
    END
END MUX4D0BWP7T

MACRO MUX4D1BWP7T
    CLASS CORE ;
    FOREIGN MUX4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.735 0.475 11.060 3.385 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.820 1.260 7.050 2.065 ;
        RECT  5.690 1.260 6.820 1.540 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.6309 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.170 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.3834 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.770 6.580 2.710 ;
        RECT  6.140 1.965 6.300 2.305 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.820 4.950 2.100 ;
        RECT  4.010 1.780 4.410 2.100 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        RECT  1.245 1.770 1.260 2.140 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2160 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 1.770 3.780 2.250 ;
        RECT  2.940 1.770 3.400 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.210 -0.235 11.200 0.235 ;
        RECT  9.870 -0.235 10.210 0.465 ;
        RECT  6.825 -0.235 9.870 0.235 ;
        RECT  6.485 -0.235 6.825 0.465 ;
        RECT  4.105 -0.235 6.485 0.235 ;
        RECT  3.765 -0.235 4.105 0.740 ;
        RECT  1.240 -0.235 3.765 0.235 ;
        RECT  0.900 -0.235 1.240 1.080 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 3.685 11.200 4.155 ;
        RECT  9.960 3.250 10.300 4.155 ;
        RECT  6.655 3.685 9.960 4.155 ;
        RECT  6.315 3.455 6.655 4.155 ;
        RECT  4.040 3.685 6.315 4.155 ;
        RECT  3.700 3.050 4.040 4.155 ;
        RECT  0.465 3.685 3.700 4.155 ;
        RECT  0.235 3.400 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.275 1.165 10.505 2.425 ;
        RECT  9.705 1.165 10.275 1.395 ;
        RECT  9.705 2.195 10.275 2.425 ;
        RECT  8.970 1.625 10.040 1.965 ;
        RECT  9.475 0.945 9.705 1.395 ;
        RECT  9.475 2.195 9.705 3.345 ;
        RECT  7.095 3.115 9.475 3.345 ;
        RECT  8.740 0.900 8.970 2.825 ;
        RECT  8.020 0.705 8.250 2.825 ;
        RECT  5.460 0.705 8.020 0.935 ;
        RECT  7.560 1.275 7.790 2.715 ;
        RECT  7.530 1.275 7.560 1.505 ;
        RECT  7.530 2.485 7.560 2.715 ;
        RECT  7.300 1.165 7.530 1.505 ;
        RECT  7.300 2.485 7.530 2.825 ;
        RECT  6.865 2.940 7.095 3.345 ;
        RECT  5.795 2.940 6.865 3.170 ;
        RECT  5.565 2.940 5.795 3.285 ;
        RECT  4.655 3.055 5.565 3.285 ;
        RECT  5.240 0.705 5.460 2.675 ;
        RECT  5.230 0.705 5.240 2.825 ;
        RECT  4.980 1.220 5.230 1.450 ;
        RECT  5.010 2.420 5.230 2.825 ;
        RECT  4.770 0.605 5.000 0.945 ;
        RECT  4.730 0.715 4.770 0.945 ;
        RECT  4.500 0.715 4.730 1.200 ;
        RECT  4.420 2.590 4.655 3.285 ;
        RECT  3.435 0.970 4.500 1.200 ;
        RECT  2.645 2.590 4.420 2.820 ;
        RECT  3.195 0.660 3.435 1.200 ;
        RECT  2.185 0.660 3.195 0.890 ;
        RECT  2.415 1.165 2.645 3.225 ;
        RECT  2.370 2.885 2.415 3.225 ;
        RECT  1.955 0.660 2.185 2.545 ;
        RECT  0.465 1.310 1.955 1.540 ;
        RECT  0.345 0.840 0.465 1.540 ;
        RECT  0.345 2.700 0.465 3.040 ;
        RECT  0.235 0.840 0.345 3.040 ;
        RECT  0.115 1.310 0.235 3.040 ;
    END
END MUX4D1BWP7T

MACRO MUX4D2BWP7T
    CLASS CORE ;
    FOREIGN MUX4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.525 1.010 17.780 2.470 ;
        RECT  17.500 0.465 17.525 3.325 ;
        RECT  17.295 0.465 17.500 1.305 ;
        RECT  17.295 2.240 17.500 3.325 ;
        END
    END Z
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.300 1.660 13.550 2.005 ;
        RECT  13.020 1.615 13.300 2.710 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.6309 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 3.225 4.465 3.455 ;
        RECT  3.035 2.985 3.275 3.455 ;
        RECT  1.375 2.985 3.035 3.225 ;
        RECT  1.095 2.480 1.375 3.225 ;
        RECT  0.980 2.480 1.095 2.710 ;
        RECT  0.700 1.635 0.980 2.710 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.615 12.740 2.150 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.8487 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.260 8.310 1.540 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.100 2.150 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.130 1.260 6.070 1.540 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 -0.235 18.480 0.235 ;
        RECT  18.015 -0.235 18.245 1.240 ;
        RECT  16.820 -0.235 18.015 0.235 ;
        RECT  16.480 -0.235 16.820 0.465 ;
        RECT  13.475 -0.235 16.480 0.235 ;
        RECT  13.095 -0.235 13.475 0.465 ;
        RECT  11.960 -0.235 13.095 0.235 ;
        RECT  11.580 -0.235 11.960 0.465 ;
        RECT  8.705 -0.235 11.580 0.235 ;
        RECT  8.365 -0.235 8.705 0.510 ;
        RECT  7.250 -0.235 8.365 0.235 ;
        RECT  6.870 -0.235 7.250 0.940 ;
        RECT  5.770 -0.235 6.870 0.235 ;
        RECT  5.390 -0.235 5.770 0.465 ;
        RECT  2.745 -0.235 5.390 0.235 ;
        RECT  2.365 -0.235 2.745 0.465 ;
        RECT  1.185 -0.235 2.365 0.235 ;
        RECT  0.955 -0.235 1.185 0.815 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 3.685 18.480 4.155 ;
        RECT  18.015 2.250 18.245 4.155 ;
        RECT  16.860 3.685 18.015 4.155 ;
        RECT  16.520 3.225 16.860 4.155 ;
        RECT  13.405 3.685 16.520 4.155 ;
        RECT  13.065 3.455 13.405 4.155 ;
        RECT  11.885 3.685 13.065 4.155 ;
        RECT  11.545 3.455 11.885 4.155 ;
        RECT  8.685 3.685 11.545 4.155 ;
        RECT  8.345 3.190 8.685 4.155 ;
        RECT  7.205 3.685 8.345 4.155 ;
        RECT  6.865 2.730 7.205 4.155 ;
        RECT  5.725 3.685 6.865 4.155 ;
        RECT  5.385 3.190 5.725 4.155 ;
        RECT  2.805 3.685 5.385 4.155 ;
        RECT  2.465 3.455 2.805 4.155 ;
        RECT  1.285 3.685 2.465 4.155 ;
        RECT  0.945 3.455 1.285 4.155 ;
        RECT  0.000 3.685 0.945 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.835 0.995 17.065 2.560 ;
        RECT  15.980 0.995 16.835 1.230 ;
        RECT  16.265 2.330 16.835 2.560 ;
        RECT  15.505 1.715 16.605 1.945 ;
        RECT  16.035 2.330 16.265 3.455 ;
        RECT  14.160 3.225 16.035 3.455 ;
        RECT  15.275 0.500 15.505 2.945 ;
        RECT  14.805 0.500 14.840 0.735 ;
        RECT  14.575 0.500 14.805 2.945 ;
        RECT  14.500 0.500 14.575 0.925 ;
        RECT  14.555 2.605 14.575 2.945 ;
        RECT  13.255 0.695 14.500 0.925 ;
        RECT  14.265 1.655 14.345 1.995 ;
        RECT  14.085 1.155 14.265 1.995 ;
        RECT  13.930 2.990 14.160 3.455 ;
        RECT  13.925 1.155 14.085 2.755 ;
        RECT  11.240 2.990 13.930 3.225 ;
        RECT  13.855 1.690 13.925 2.755 ;
        RECT  13.025 0.695 13.255 1.385 ;
        RECT  10.430 1.155 13.025 1.385 ;
        RECT  10.745 2.530 12.645 2.760 ;
        RECT  12.405 0.500 12.635 0.925 ;
        RECT  10.865 0.695 12.405 0.925 ;
        RECT  10.960 2.990 11.240 3.300 ;
        RECT  9.850 3.045 10.960 3.300 ;
        RECT  10.310 0.700 10.430 2.705 ;
        RECT  10.200 0.700 10.310 2.815 ;
        RECT  10.080 2.475 10.200 2.815 ;
        RECT  9.620 2.270 9.850 3.300 ;
        RECT  9.420 1.400 9.650 2.030 ;
        RECT  4.225 2.270 9.620 2.500 ;
        RECT  7.605 0.740 9.465 0.970 ;
        RECT  4.690 1.800 9.420 2.030 ;
        RECT  9.160 2.730 9.390 3.070 ;
        RECT  7.585 2.730 9.160 2.960 ;
        RECT  4.645 0.755 6.505 0.985 ;
        RECT  4.625 2.730 6.485 2.960 ;
        RECT  4.460 1.415 4.690 2.030 ;
        RECT  4.170 2.270 4.225 2.780 ;
        RECT  3.940 0.965 4.170 2.780 ;
        RECT  3.885 2.490 3.940 2.780 ;
        RECT  3.215 0.695 3.445 1.330 ;
        RECT  1.705 2.490 3.340 2.720 ;
        RECT  1.905 0.695 3.215 0.925 ;
        RECT  2.595 1.620 3.010 1.850 ;
        RECT  2.365 1.155 2.595 1.850 ;
        RECT  0.465 1.155 2.365 1.385 ;
        RECT  1.675 0.510 1.905 0.925 ;
        RECT  0.235 0.475 0.465 3.025 ;
    END
END MUX4D2BWP7T

MACRO MUX4ND0BWP7T
    CLASS CORE ;
    FOREIGN MUX4ND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6552 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.110 1.210 9.380 2.710 ;
        RECT  9.100 0.900 9.110 2.825 ;
        RECT  8.880 0.900 9.100 1.440 ;
        RECT  8.880 2.480 9.100 2.825 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.960 1.260 7.190 2.065 ;
        RECT  6.250 1.260 6.960 1.540 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.6399 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.170 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.3303 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.770 6.580 2.710 ;
        RECT  6.280 1.965 6.300 2.305 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.2673 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.365 1.820 5.250 2.100 ;
        RECT  4.010 1.780 4.365 2.100 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.2655 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        RECT  1.245 1.770 1.260 2.140 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 1.770 3.780 2.150 ;
        RECT  3.355 1.770 3.695 2.265 ;
        RECT  2.940 1.770 3.355 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.965 -0.235 10.080 0.235 ;
        RECT  6.625 -0.235 6.965 0.465 ;
        RECT  4.105 -0.235 6.625 0.235 ;
        RECT  3.765 -0.235 4.105 0.740 ;
        RECT  1.240 -0.235 3.765 0.235 ;
        RECT  0.900 -0.235 1.240 1.080 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.785 3.685 10.080 4.155 ;
        RECT  6.555 3.400 6.785 4.155 ;
        RECT  3.975 3.685 6.555 4.155 ;
        RECT  3.635 3.050 3.975 4.155 ;
        RECT  1.240 3.685 3.635 4.155 ;
        RECT  0.900 3.250 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.615 0.870 9.845 3.345 ;
        RECT  7.240 3.115 9.615 3.345 ;
        RECT  8.160 0.705 8.390 2.825 ;
        RECT  5.760 0.705 8.160 0.935 ;
        RECT  7.700 1.275 7.930 2.715 ;
        RECT  7.670 1.275 7.700 1.505 ;
        RECT  7.670 2.485 7.700 2.715 ;
        RECT  7.440 1.165 7.670 1.505 ;
        RECT  7.440 2.485 7.670 2.825 ;
        RECT  7.010 2.940 7.240 3.345 ;
        RECT  5.855 2.940 7.010 3.170 ;
        RECT  5.625 2.940 5.855 3.285 ;
        RECT  5.530 0.705 5.760 2.675 ;
        RECT  4.930 3.055 5.625 3.285 ;
        RECT  5.335 1.220 5.530 1.450 ;
        RECT  5.410 2.420 5.530 2.675 ;
        RECT  5.180 2.420 5.410 2.825 ;
        RECT  5.070 0.605 5.300 0.945 ;
        RECT  4.570 0.715 5.070 0.945 ;
        RECT  4.695 2.590 4.930 3.285 ;
        RECT  2.635 2.590 4.695 2.820 ;
        RECT  4.340 0.715 4.570 1.200 ;
        RECT  3.145 0.970 4.340 1.200 ;
        RECT  2.905 0.660 3.145 1.200 ;
        RECT  2.000 0.660 2.905 0.890 ;
        RECT  2.405 1.165 2.635 3.225 ;
        RECT  2.230 2.885 2.405 3.225 ;
        RECT  2.000 2.205 2.145 2.545 ;
        RECT  1.770 0.660 2.000 2.545 ;
        RECT  0.465 1.310 1.770 1.540 ;
        RECT  0.345 3.110 0.520 3.340 ;
        RECT  0.345 0.840 0.465 1.540 ;
        RECT  0.235 0.840 0.345 3.340 ;
        RECT  0.115 1.310 0.235 3.340 ;
    END
END MUX4ND0BWP7T

MACRO MUX4ND1BWP7T
    CLASS CORE ;
    FOREIGN MUX4ND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.975 0.475 13.300 3.385 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.770 9.380 2.150 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.6309 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.170 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.3834 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.770 6.580 2.710 ;
        RECT  6.020 1.885 6.300 2.225 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.820 4.950 2.100 ;
        RECT  4.010 1.780 4.410 2.100 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        RECT  1.245 1.770 1.260 2.140 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 1.770 3.780 2.250 ;
        RECT  2.940 1.770 3.400 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.450 -0.235 13.440 0.235 ;
        RECT  12.110 -0.235 12.450 0.465 ;
        RECT  9.065 -0.235 12.110 0.235 ;
        RECT  8.725 -0.235 9.065 0.465 ;
        RECT  6.825 -0.235 8.725 0.235 ;
        RECT  6.485 -0.235 6.825 0.465 ;
        RECT  4.105 -0.235 6.485 0.235 ;
        RECT  3.765 -0.235 4.105 0.740 ;
        RECT  1.240 -0.235 3.765 0.235 ;
        RECT  0.900 -0.235 1.240 1.080 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.540 3.685 13.440 4.155 ;
        RECT  12.200 3.250 12.540 4.155 ;
        RECT  9.065 3.685 12.200 4.155 ;
        RECT  8.725 3.455 9.065 4.155 ;
        RECT  6.655 3.685 8.725 4.155 ;
        RECT  6.315 3.455 6.655 4.155 ;
        RECT  4.040 3.685 6.315 4.155 ;
        RECT  3.700 3.050 4.040 4.155 ;
        RECT  0.465 3.685 3.700 4.155 ;
        RECT  0.235 3.400 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.515 1.165 12.745 2.425 ;
        RECT  11.945 1.165 12.515 1.395 ;
        RECT  11.945 2.195 12.515 2.425 ;
        RECT  11.225 1.625 12.280 1.965 ;
        RECT  11.715 0.945 11.945 1.395 ;
        RECT  11.715 2.195 11.945 3.375 ;
        RECT  9.750 3.145 11.715 3.375 ;
        RECT  10.995 0.900 11.225 2.825 ;
        RECT  10.275 0.695 10.505 2.825 ;
        RECT  7.530 0.695 10.275 0.925 ;
        RECT  9.805 1.155 10.030 2.610 ;
        RECT  9.800 1.155 9.805 2.720 ;
        RECT  9.520 1.155 9.800 1.385 ;
        RECT  9.575 2.380 9.800 2.720 ;
        RECT  9.500 2.995 9.750 3.375 ;
        RECT  8.195 2.995 9.500 3.225 ;
        RECT  8.195 1.155 8.305 1.385 ;
        RECT  7.965 1.155 8.195 3.225 ;
        RECT  7.500 2.995 7.730 3.430 ;
        RECT  7.300 0.695 7.530 2.755 ;
        RECT  5.795 2.995 7.500 3.225 ;
        RECT  7.075 2.525 7.300 2.755 ;
        RECT  6.820 1.220 7.050 2.065 ;
        RECT  5.460 1.220 6.820 1.450 ;
        RECT  5.565 2.995 5.795 3.285 ;
        RECT  4.655 3.055 5.565 3.285 ;
        RECT  5.240 1.220 5.460 2.675 ;
        RECT  5.230 1.220 5.240 2.825 ;
        RECT  4.980 1.220 5.230 1.450 ;
        RECT  5.010 2.420 5.230 2.825 ;
        RECT  4.770 0.605 5.000 0.945 ;
        RECT  4.730 0.715 4.770 0.945 ;
        RECT  4.500 0.715 4.730 1.200 ;
        RECT  4.420 2.590 4.655 3.285 ;
        RECT  3.435 0.970 4.500 1.200 ;
        RECT  2.645 2.590 4.420 2.820 ;
        RECT  3.195 0.660 3.435 1.200 ;
        RECT  2.185 0.660 3.195 0.890 ;
        RECT  2.415 1.165 2.645 3.225 ;
        RECT  2.370 2.885 2.415 3.225 ;
        RECT  1.955 0.660 2.185 2.545 ;
        RECT  0.465 1.310 1.955 1.540 ;
        RECT  0.345 0.840 0.465 1.540 ;
        RECT  0.345 2.700 0.465 3.040 ;
        RECT  0.235 0.840 0.345 3.040 ;
        RECT  0.115 1.310 0.235 3.040 ;
    END
END MUX4ND1BWP7T

MACRO MUX4ND2BWP7T
    CLASS CORE ;
    FOREIGN MUX4ND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.045 1.210 13.300 2.150 ;
        RECT  12.815 0.475 13.045 3.385 ;
        END
    END ZN
    PIN S1
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.770 9.380 2.150 ;
        END
    END S1
    PIN S0
        ANTENNAGATEAREA 0.6309 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.575 1.770 0.700 2.170 ;
        END
    END S0
    PIN I3
        ANTENNAGATEAREA 0.3834 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.770 6.580 2.710 ;
        RECT  6.020 1.885 6.300 2.225 ;
        END
    END I3
    PIN I2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.820 4.950 2.100 ;
        RECT  4.010 1.780 4.410 2.100 ;
        END
    END I2
    PIN I1
        ANTENNAGATEAREA 0.3456 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        RECT  1.245 1.770 1.260 2.140 ;
        END
    END I1
    PIN I0
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 1.770 3.780 2.250 ;
        RECT  2.940 1.770 3.400 2.150 ;
        END
    END I0
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.765 -0.235 14.000 0.235 ;
        RECT  13.535 -0.235 13.765 1.285 ;
        RECT  12.290 -0.235 13.535 0.235 ;
        RECT  11.950 -0.235 12.290 0.465 ;
        RECT  9.045 -0.235 11.950 0.235 ;
        RECT  8.705 -0.235 9.045 0.465 ;
        RECT  6.825 -0.235 8.705 0.235 ;
        RECT  6.485 -0.235 6.825 0.465 ;
        RECT  4.105 -0.235 6.485 0.235 ;
        RECT  3.765 -0.235 4.105 0.740 ;
        RECT  1.240 -0.235 3.765 0.235 ;
        RECT  0.900 -0.235 1.240 1.080 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.765 3.685 14.000 4.155 ;
        RECT  13.535 2.255 13.765 4.155 ;
        RECT  12.380 3.685 13.535 4.155 ;
        RECT  12.040 3.250 12.380 4.155 ;
        RECT  8.975 3.685 12.040 4.155 ;
        RECT  8.635 3.455 8.975 4.155 ;
        RECT  6.655 3.685 8.635 4.155 ;
        RECT  6.315 3.455 6.655 4.155 ;
        RECT  4.040 3.685 6.315 4.155 ;
        RECT  3.700 3.050 4.040 4.155 ;
        RECT  0.465 3.685 3.700 4.155 ;
        RECT  0.235 3.400 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.355 1.165 12.585 2.425 ;
        RECT  11.785 1.165 12.355 1.395 ;
        RECT  11.785 2.195 12.355 2.425 ;
        RECT  11.065 1.625 12.120 1.965 ;
        RECT  11.555 0.945 11.785 1.395 ;
        RECT  11.555 2.195 11.785 3.375 ;
        RECT  9.590 3.145 11.555 3.375 ;
        RECT  10.835 0.900 11.065 2.825 ;
        RECT  10.115 0.695 10.345 2.825 ;
        RECT  7.530 0.695 10.115 0.925 ;
        RECT  9.645 1.155 9.870 2.610 ;
        RECT  9.640 1.155 9.645 2.720 ;
        RECT  9.360 1.155 9.640 1.385 ;
        RECT  9.415 2.380 9.640 2.720 ;
        RECT  9.340 2.995 9.590 3.375 ;
        RECT  9.065 2.995 9.340 3.225 ;
        RECT  8.835 2.565 9.065 3.225 ;
        RECT  8.160 2.565 8.835 2.795 ;
        RECT  8.160 1.155 8.285 1.385 ;
        RECT  7.930 1.155 8.160 2.795 ;
        RECT  7.490 2.995 7.720 3.430 ;
        RECT  7.300 0.695 7.530 2.755 ;
        RECT  5.795 2.995 7.490 3.225 ;
        RECT  7.075 2.525 7.300 2.755 ;
        RECT  6.820 1.220 7.050 2.065 ;
        RECT  5.460 1.220 6.820 1.450 ;
        RECT  5.565 2.995 5.795 3.285 ;
        RECT  4.655 3.055 5.565 3.285 ;
        RECT  5.240 1.220 5.460 2.675 ;
        RECT  5.230 1.220 5.240 2.825 ;
        RECT  4.980 1.220 5.230 1.450 ;
        RECT  5.010 2.420 5.230 2.825 ;
        RECT  4.770 0.605 5.000 0.945 ;
        RECT  4.730 0.715 4.770 0.945 ;
        RECT  4.500 0.715 4.730 1.200 ;
        RECT  4.420 2.590 4.655 3.285 ;
        RECT  3.435 0.970 4.500 1.200 ;
        RECT  2.645 2.590 4.420 2.820 ;
        RECT  3.195 0.660 3.435 1.200 ;
        RECT  2.185 0.660 3.195 0.890 ;
        RECT  2.415 1.165 2.645 3.225 ;
        RECT  2.370 2.885 2.415 3.225 ;
        RECT  1.955 0.660 2.185 2.545 ;
        RECT  0.465 1.310 1.955 1.540 ;
        RECT  0.345 2.700 0.465 3.040 ;
        RECT  0.235 0.840 0.345 3.040 ;
        RECT  0.115 1.310 0.235 3.040 ;
        RECT  0.345 0.840 0.465 1.540 ;
    END
END MUX4ND2BWP7T

MACRO ND2D0BWP7T
    CLASS CORE ;
    FOREIGN ND2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6099 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 0.580 1.920 0.810 ;
        RECT  1.260 0.580 1.540 2.150 ;
        RECT  1.225 1.820 1.260 2.150 ;
        RECT  0.995 1.820 1.225 3.145 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 1.210 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 -0.235 2.240 0.235 ;
        RECT  0.270 -0.235 0.510 0.865 ;
        RECT  0.000 -0.235 0.270 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 3.685 2.240 4.155 ;
        RECT  1.710 2.800 1.950 4.155 ;
        RECT  0.510 3.685 1.710 4.155 ;
        RECT  0.270 2.805 0.510 4.155 ;
        RECT  0.000 3.685 0.270 4.155 ;
        END
    END VDD
END ND2D0BWP7T

MACRO ND2D1BWP7T
    CLASS CORE ;
    FOREIGN ND2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2198 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 0.750 1.920 0.980 ;
        RECT  1.260 0.750 1.540 2.150 ;
        RECT  1.225 1.820 1.260 2.150 ;
        RECT  0.995 1.820 1.225 3.385 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 1.210 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 -0.235 2.240 0.235 ;
        RECT  0.270 -0.235 0.510 0.930 ;
        RECT  0.000 -0.235 0.270 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 3.685 2.240 4.155 ;
        RECT  1.710 2.510 1.950 4.155 ;
        RECT  0.510 3.685 1.710 4.155 ;
        RECT  0.270 2.470 0.510 4.155 ;
        RECT  0.000 3.685 0.270 4.155 ;
        END
    END VDD
END ND2D1BWP7T

MACRO ND2D1P5BWP7T
    CLASS CORE ;
    FOREIGN ND2D1P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.5147 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 2.380 2.880 2.610 ;
        RECT  1.925 0.770 2.100 2.610 ;
        RECT  1.820 0.565 1.925 2.610 ;
        RECT  1.695 0.565 1.820 0.975 ;
        RECT  1.020 2.380 1.820 2.610 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.6399 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.140 1.715 3.380 3.070 ;
        RECT  2.730 1.715 3.140 1.945 ;
        RECT  0.455 2.840 3.140 3.070 ;
        RECT  0.140 1.210 0.455 3.070 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6399 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.715 1.590 1.945 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.330 -0.235 3.920 0.235 ;
        RECT  2.950 -0.235 3.330 0.770 ;
        RECT  0.660 -0.235 2.950 0.235 ;
        RECT  0.280 -0.235 0.660 0.770 ;
        RECT  0.000 -0.235 0.280 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.740 3.685 3.920 4.155 ;
        RECT  3.400 3.300 3.740 4.155 ;
        RECT  2.120 3.685 3.400 4.155 ;
        RECT  1.780 3.300 2.120 4.155 ;
        RECT  0.520 3.685 1.780 4.155 ;
        RECT  0.180 3.300 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
END ND2D1P5BWP7T

MACRO ND2D2BWP7T
    CLASS CORE ;
    FOREIGN ND2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.1396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 2.300 2.880 2.530 ;
        RECT  2.380 1.020 2.660 2.530 ;
        RECT  2.045 1.020 2.380 1.250 ;
        RECT  0.980 2.300 2.380 2.530 ;
        RECT  1.815 0.635 2.045 1.250 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.235 1.585 3.465 2.990 ;
        RECT  0.455 2.760 3.235 2.990 ;
        RECT  0.140 1.585 0.455 2.990 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.640 1.990 1.870 ;
        RECT  1.260 0.650 1.540 1.870 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.640 -0.235 3.920 0.235 ;
        RECT  3.260 -0.235 3.640 1.195 ;
        RECT  0.580 -0.235 3.260 0.235 ;
        RECT  0.200 -0.235 0.580 1.195 ;
        RECT  0.000 -0.235 0.200 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.660 3.685 3.920 4.155 ;
        RECT  3.315 3.220 3.660 4.155 ;
        RECT  2.100 3.685 3.315 4.155 ;
        RECT  1.720 3.220 2.100 4.155 ;
        RECT  0.560 3.685 1.720 4.155 ;
        RECT  0.220 3.220 0.560 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
END ND2D2BWP7T

MACRO ND2D2P5BWP7T
    CLASS CORE ;
    FOREIGN ND2D2P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.7179 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 0.750 4.900 2.800 ;
        RECT  2.670 0.750 4.575 0.980 ;
        RECT  4.065 2.560 4.575 2.800 ;
        RECT  3.835 2.560 4.065 3.455 ;
        RECT  2.625 2.560 3.835 2.800 ;
        RECT  2.440 0.585 2.670 0.980 ;
        RECT  2.395 2.560 2.625 3.440 ;
        RECT  1.660 0.585 2.440 0.815 ;
        RECT  0.890 2.560 2.395 2.790 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.0674 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.140 1.620 3.625 1.850 ;
        RECT  1.910 1.125 2.140 1.850 ;
        RECT  0.470 1.125 1.910 1.355 ;
        RECT  0.140 1.125 0.470 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.0674 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.330 ;
        RECT  1.540 2.080 4.060 2.330 ;
        RECT  1.260 1.585 1.540 2.330 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.480 -0.235 5.040 0.235 ;
        RECT  3.020 -0.235 3.480 0.520 ;
        RECT  0.580 -0.235 3.020 0.235 ;
        RECT  0.200 -0.235 0.580 0.845 ;
        RECT  0.000 -0.235 0.200 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 3.685 5.040 4.155 ;
        RECT  4.500 3.115 4.880 4.155 ;
        RECT  3.440 3.685 4.500 4.155 ;
        RECT  3.060 3.110 3.440 4.155 ;
        RECT  1.960 3.685 3.060 4.155 ;
        RECT  1.620 3.100 1.960 4.155 ;
        RECT  0.465 3.685 1.620 4.155 ;
        RECT  0.235 2.525 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
END ND2D2P5BWP7T

MACRO ND2D3BWP7T
    CLASS CORE ;
    FOREIGN ND2D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.2394 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.555 0.495 4.785 1.375 ;
        RECT  4.065 1.015 4.555 1.375 ;
        RECT  3.835 1.015 4.065 3.330 ;
        RECT  3.190 1.015 3.835 2.780 ;
        RECT  3.060 1.015 3.190 1.365 ;
        RECT  2.625 2.430 3.190 2.780 ;
        RECT  2.395 2.430 2.625 3.330 ;
        RECT  1.185 2.430 2.395 2.780 ;
        RECT  0.955 2.430 1.185 3.330 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.655 1.735 2.220 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.715 4.900 2.710 ;
        RECT  4.370 1.715 4.620 1.945 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 -0.235 5.040 0.235 ;
        RECT  1.605 -0.235 1.985 0.785 ;
        RECT  0.560 -0.235 1.605 0.235 ;
        RECT  0.180 -0.235 0.560 1.250 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.865 3.685 5.040 4.155 ;
        RECT  4.485 3.045 4.865 4.155 ;
        RECT  3.435 3.685 4.485 4.155 ;
        RECT  3.055 3.045 3.435 4.155 ;
        RECT  1.995 3.685 3.055 4.155 ;
        RECT  1.615 3.045 1.995 4.155 ;
        RECT  0.555 3.685 1.615 4.155 ;
        RECT  0.175 2.485 0.555 4.155 ;
        RECT  0.000 3.685 0.175 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.625 0.495 4.120 0.725 ;
        RECT  2.395 0.495 2.625 1.305 ;
        RECT  1.185 1.035 2.395 1.305 ;
        RECT  0.955 0.495 1.185 1.305 ;
    END
END ND2D3BWP7T

MACRO ND2D4BWP7T
    CLASS CORE ;
    FOREIGN ND2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 4.0511 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.650 1.020 5.665 1.250 ;
        RECT  5.380 2.380 5.610 3.240 ;
        RECT  4.650 2.380 5.380 2.730 ;
        RECT  4.170 1.020 4.650 2.730 ;
        RECT  3.940 1.020 4.170 3.240 ;
        RECT  3.750 1.020 3.940 2.730 ;
        RECT  2.725 2.380 3.750 2.730 ;
        RECT  2.495 2.380 2.725 3.240 ;
        RECT  1.285 2.380 2.495 2.730 ;
        RECT  1.055 2.380 1.285 3.240 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.625 2.855 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.060 1.625 6.020 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.810 -0.235 6.720 0.235 ;
        RECT  2.430 -0.235 2.810 0.810 ;
        RECT  1.370 -0.235 2.430 0.235 ;
        RECT  0.990 -0.235 1.370 0.810 ;
        RECT  0.000 -0.235 0.990 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.420 3.685 6.720 4.155 ;
        RECT  6.040 2.485 6.420 4.155 ;
        RECT  4.980 3.685 6.040 4.155 ;
        RECT  4.600 2.960 4.980 4.155 ;
        RECT  3.540 3.685 4.600 4.155 ;
        RECT  3.160 2.960 3.540 4.155 ;
        RECT  2.100 3.685 3.160 4.155 ;
        RECT  1.720 2.960 2.100 4.155 ;
        RECT  0.660 3.685 1.720 4.155 ;
        RECT  0.280 2.485 0.660 4.155 ;
        RECT  0.000 3.685 0.280 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.850 1.020 5.665 1.250 ;
        RECT  5.380 2.380 5.610 3.240 ;
        RECT  4.850 2.380 5.380 2.730 ;
        RECT  2.725 2.380 3.550 2.730 ;
        RECT  2.495 2.380 2.725 3.240 ;
        RECT  1.285 2.380 2.495 2.730 ;
        RECT  1.055 2.380 1.285 3.240 ;
        RECT  6.100 0.475 6.330 1.285 ;
        RECT  3.445 0.475 6.100 0.715 ;
        RECT  3.215 0.475 3.445 1.300 ;
        RECT  2.065 1.070 3.215 1.300 ;
        RECT  1.720 0.540 2.065 1.300 ;
        RECT  0.625 1.070 1.720 1.300 ;
        RECT  0.280 0.500 0.625 1.300 ;
    END
END ND2D4BWP7T

MACRO ND2D5BWP7T
    CLASS CORE ;
    FOREIGN ND2D5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.2640 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.590 0.495 7.955 1.345 ;
        RECT  5.770 1.020 7.590 1.345 ;
        RECT  6.940 2.400 7.170 3.295 ;
        RECT  5.770 2.400 6.940 2.750 ;
        RECT  5.730 1.020 5.770 2.750 ;
        RECT  5.500 1.020 5.730 3.295 ;
        RECT  4.870 1.020 5.500 2.750 ;
        RECT  4.670 1.020 4.870 1.345 ;
        RECT  4.285 2.400 4.870 2.750 ;
        RECT  4.055 2.400 4.285 3.295 ;
        RECT  2.845 2.400 4.055 2.750 ;
        RECT  2.615 2.400 2.845 3.295 ;
        RECT  1.405 2.400 2.615 2.750 ;
        RECT  1.175 2.400 1.405 3.295 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 2.1330 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 1.610 3.575 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.1330 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.140 1.610 7.410 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.650 -0.235 8.400 0.235 ;
        RECT  3.270 -0.235 3.650 0.785 ;
        RECT  2.210 -0.235 3.270 0.235 ;
        RECT  1.830 -0.235 2.210 0.785 ;
        RECT  0.760 -0.235 1.830 0.235 ;
        RECT  0.380 -0.235 0.760 1.195 ;
        RECT  0.000 -0.235 0.380 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 3.685 8.400 4.155 ;
        RECT  7.600 2.540 7.980 4.155 ;
        RECT  6.540 3.685 7.600 4.155 ;
        RECT  6.160 2.980 6.540 4.155 ;
        RECT  5.100 3.685 6.160 4.155 ;
        RECT  4.720 2.980 5.100 4.155 ;
        RECT  3.660 3.685 4.720 4.155 ;
        RECT  3.280 2.980 3.660 4.155 ;
        RECT  2.220 3.685 3.280 4.155 ;
        RECT  1.840 2.980 2.220 4.155 ;
        RECT  0.780 3.685 1.840 4.155 ;
        RECT  0.400 2.540 0.780 4.155 ;
        RECT  0.000 3.685 0.400 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.590 0.495 7.955 1.345 ;
        RECT  5.970 1.020 7.590 1.345 ;
        RECT  6.940 2.400 7.170 3.295 ;
        RECT  5.970 2.400 6.940 2.750 ;
        RECT  4.285 2.400 4.670 2.750 ;
        RECT  4.055 2.400 4.285 3.295 ;
        RECT  2.845 2.400 4.055 2.750 ;
        RECT  2.615 2.400 2.845 3.295 ;
        RECT  1.405 2.400 2.615 2.750 ;
        RECT  1.175 2.400 1.405 3.295 ;
        RECT  4.285 0.465 7.225 0.695 ;
        RECT  4.055 0.465 4.285 1.310 ;
        RECT  2.900 1.040 4.055 1.310 ;
        RECT  2.560 0.490 2.900 1.310 ;
        RECT  1.460 1.040 2.560 1.310 ;
        RECT  1.120 0.495 1.460 1.310 ;
    END
END ND2D5BWP7T

MACRO ND2D6BWP7T
    CLASS CORE ;
    FOREIGN ND2D6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 6.0706 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.330 0.965 8.410 1.315 ;
        RECT  8.180 2.400 8.410 3.330 ;
        RECT  6.970 2.400 8.180 2.750 ;
        RECT  6.740 2.400 6.970 3.330 ;
        RECT  6.330 2.400 6.740 2.750 ;
        RECT  5.530 0.965 6.330 2.750 ;
        RECT  5.430 0.965 5.530 3.330 ;
        RECT  5.245 0.965 5.430 1.315 ;
        RECT  5.300 2.400 5.430 3.330 ;
        RECT  4.085 2.400 5.300 2.750 ;
        RECT  3.855 2.400 4.085 3.330 ;
        RECT  2.645 2.400 3.855 2.750 ;
        RECT  2.415 2.400 2.645 3.330 ;
        RECT  1.205 2.400 2.415 2.750 ;
        RECT  0.975 2.400 1.205 3.330 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 2.5596 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.735 1.655 4.255 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.5596 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.770 1.655 8.410 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.170 -0.235 9.520 0.235 ;
        RECT  3.790 -0.235 4.170 0.785 ;
        RECT  2.730 -0.235 3.790 0.235 ;
        RECT  2.350 -0.235 2.730 0.785 ;
        RECT  1.290 -0.235 2.350 0.235 ;
        RECT  0.910 -0.235 1.290 0.785 ;
        RECT  0.000 -0.235 0.910 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.225 3.685 9.520 4.155 ;
        RECT  8.840 2.485 9.225 4.155 ;
        RECT  7.785 3.685 8.840 4.155 ;
        RECT  7.400 3.045 7.785 4.155 ;
        RECT  6.345 3.685 7.400 4.155 ;
        RECT  5.960 3.045 6.345 4.155 ;
        RECT  4.900 3.685 5.960 4.155 ;
        RECT  4.515 3.045 4.900 4.155 ;
        RECT  3.460 3.685 4.515 4.155 ;
        RECT  3.075 3.045 3.460 4.155 ;
        RECT  2.020 3.685 3.075 4.155 ;
        RECT  1.635 3.045 2.020 4.155 ;
        RECT  0.580 3.685 1.635 4.155 ;
        RECT  0.200 2.450 0.580 4.155 ;
        RECT  0.000 3.685 0.200 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.530 0.965 8.410 1.315 ;
        RECT  8.180 2.400 8.410 3.330 ;
        RECT  6.970 2.400 8.180 2.750 ;
        RECT  6.740 2.400 6.970 3.330 ;
        RECT  6.530 2.400 6.740 2.750 ;
        RECT  4.085 2.400 5.230 2.750 ;
        RECT  3.855 2.400 4.085 3.330 ;
        RECT  2.645 2.400 3.855 2.750 ;
        RECT  2.415 2.400 2.645 3.330 ;
        RECT  1.205 2.400 2.415 2.750 ;
        RECT  0.975 2.400 1.205 3.330 ;
        RECT  8.900 0.465 9.130 1.275 ;
        RECT  4.805 0.465 8.900 0.725 ;
        RECT  4.575 0.465 4.805 1.360 ;
        RECT  3.420 1.040 4.575 1.360 ;
        RECT  3.080 0.495 3.420 1.360 ;
        RECT  1.980 1.040 3.080 1.360 ;
        RECT  1.640 0.495 1.980 1.360 ;
        RECT  0.540 1.040 1.640 1.360 ;
        RECT  0.200 0.495 0.540 1.360 ;
    END
END ND2D6BWP7T

MACRO ND2D8BWP7T
    CLASS CORE ;
    FOREIGN ND2D8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 8.0902 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.450 0.965 11.290 1.315 ;
        RECT  11.060 2.430 11.290 3.265 ;
        RECT  9.850 2.430 11.060 2.780 ;
        RECT  9.620 2.430 9.850 3.265 ;
        RECT  8.410 2.430 9.620 2.780 ;
        RECT  8.180 2.430 8.410 3.265 ;
        RECT  7.450 2.430 8.180 2.780 ;
        RECT  6.970 0.965 7.450 2.780 ;
        RECT  6.740 0.965 6.970 3.270 ;
        RECT  6.550 0.965 6.740 2.780 ;
        RECT  5.525 2.430 6.550 2.780 ;
        RECT  5.295 2.430 5.525 3.265 ;
        RECT  4.085 2.430 5.295 2.780 ;
        RECT  3.855 2.430 4.085 3.265 ;
        RECT  2.645 2.430 3.855 2.780 ;
        RECT  2.415 2.430 2.645 3.265 ;
        RECT  1.205 2.430 2.415 2.780 ;
        RECT  0.975 2.430 1.205 3.265 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 3.4128 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.790 1.605 5.720 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 3.4128 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.880 1.610 11.400 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.610 -0.235 12.320 0.235 ;
        RECT  5.230 -0.235 5.610 0.785 ;
        RECT  4.170 -0.235 5.230 0.235 ;
        RECT  3.790 -0.235 4.170 0.785 ;
        RECT  2.730 -0.235 3.790 0.235 ;
        RECT  2.350 -0.235 2.730 0.785 ;
        RECT  1.290 -0.235 2.350 0.235 ;
        RECT  0.910 -0.235 1.290 0.785 ;
        RECT  0.000 -0.235 0.910 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.105 3.685 12.320 4.155 ;
        RECT  11.720 2.300 12.105 4.155 ;
        RECT  10.665 3.685 11.720 4.155 ;
        RECT  10.280 3.045 10.665 4.155 ;
        RECT  9.225 3.685 10.280 4.155 ;
        RECT  8.840 3.045 9.225 4.155 ;
        RECT  7.785 3.685 8.840 4.155 ;
        RECT  7.400 3.045 7.785 4.155 ;
        RECT  6.340 3.685 7.400 4.155 ;
        RECT  5.955 3.045 6.340 4.155 ;
        RECT  4.900 3.685 5.955 4.155 ;
        RECT  4.515 3.045 4.900 4.155 ;
        RECT  3.460 3.685 4.515 4.155 ;
        RECT  3.075 3.045 3.460 4.155 ;
        RECT  2.020 3.685 3.075 4.155 ;
        RECT  1.635 3.045 2.020 4.155 ;
        RECT  0.580 3.685 1.635 4.155 ;
        RECT  0.195 2.300 0.580 4.155 ;
        RECT  0.000 3.685 0.195 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.650 0.965 11.290 1.315 ;
        RECT  11.060 2.430 11.290 3.265 ;
        RECT  9.850 2.430 11.060 2.780 ;
        RECT  9.620 2.430 9.850 3.265 ;
        RECT  8.410 2.430 9.620 2.780 ;
        RECT  8.180 2.430 8.410 3.265 ;
        RECT  7.650 2.430 8.180 2.780 ;
        RECT  5.525 2.430 6.350 2.780 ;
        RECT  5.295 2.430 5.525 3.265 ;
        RECT  4.085 2.430 5.295 2.780 ;
        RECT  3.855 2.430 4.085 3.265 ;
        RECT  2.645 2.430 3.855 2.780 ;
        RECT  2.415 2.430 2.645 3.265 ;
        RECT  1.205 2.430 2.415 2.780 ;
        RECT  0.975 2.430 1.205 3.265 ;
        RECT  11.780 0.465 12.010 1.275 ;
        RECT  6.245 0.465 11.780 0.720 ;
        RECT  6.015 0.465 6.245 1.360 ;
        RECT  4.860 1.040 6.015 1.360 ;
        RECT  4.520 0.490 4.860 1.360 ;
        RECT  3.420 1.040 4.520 1.360 ;
        RECT  3.080 0.495 3.420 1.360 ;
        RECT  1.980 1.040 3.080 1.360 ;
        RECT  1.640 0.495 1.980 1.360 ;
        RECT  0.540 1.040 1.640 1.360 ;
        RECT  0.200 0.495 0.540 1.360 ;
    END
END ND2D8BWP7T

MACRO ND3D0BWP7T
    CLASS CORE ;
    FOREIGN ND3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9412 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 0.625 2.660 3.205 ;
        RECT  2.155 0.625 2.335 0.855 ;
        RECT  0.900 2.975 2.335 3.205 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 0.650 1.540 1.590 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.520 -0.235 2.800 0.235 ;
        RECT  0.180 -0.235 0.520 0.855 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 3.685 2.800 4.155 ;
        RECT  1.640 3.455 2.005 4.155 ;
        RECT  0.540 3.685 1.640 4.155 ;
        RECT  0.160 3.015 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
END ND3D0BWP7T

MACRO ND3D1BWP7T
    CLASS CORE ;
    FOREIGN ND3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.0046 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.120 3.220 2.710 ;
        RECT  2.560 1.120 2.940 1.400 ;
        RECT  2.765 2.430 2.940 2.710 ;
        RECT  2.525 2.430 2.765 3.350 ;
        RECT  2.330 0.495 2.560 1.400 ;
        RECT  1.315 2.430 2.525 2.710 ;
        RECT  1.085 2.430 1.315 3.350 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.715 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.690 -0.235 3.360 0.235 ;
        RECT  0.310 -0.235 0.690 1.190 ;
        RECT  0.000 -0.235 0.310 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 3.685 3.360 4.155 ;
        RECT  1.740 3.015 2.120 4.155 ;
        RECT  0.650 3.685 1.740 4.155 ;
        RECT  0.310 2.470 0.650 4.155 ;
        RECT  0.000 3.685 0.310 4.155 ;
        END
    END VDD
END ND3D1BWP7T

MACRO ND3D2BWP7T
    CLASS CORE ;
    FOREIGN ND3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.8394 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.065 1.320 4.340 3.020 ;
        RECT  4.060 1.320 4.065 3.445 ;
        RECT  3.630 1.320 4.060 1.550 ;
        RECT  3.835 2.790 4.060 3.445 ;
        RECT  2.625 2.790 3.835 3.020 ;
        RECT  3.400 0.925 3.630 1.550 ;
        RECT  2.340 0.925 3.400 1.155 ;
        RECT  2.395 2.790 2.625 3.445 ;
        RECT  1.185 2.790 2.395 3.020 ;
        RECT  0.955 2.790 1.185 3.445 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.570 0.860 4.800 2.000 ;
        RECT  4.125 0.860 4.570 1.090 ;
        RECT  3.895 0.465 4.125 1.090 ;
        RECT  0.980 0.465 3.895 0.695 ;
        RECT  0.700 0.465 0.980 2.150 ;
        RECT  0.640 1.530 0.700 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.480 1.780 3.590 2.010 ;
        RECT  3.250 1.780 3.480 2.560 ;
        RECT  1.540 2.330 3.250 2.560 ;
        RECT  1.260 1.155 1.540 2.560 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.770 2.710 2.100 ;
        RECT  1.820 1.210 2.100 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 -0.235 5.040 0.235 ;
        RECT  4.440 -0.235 4.880 0.630 ;
        RECT  0.465 -0.235 4.440 0.235 ;
        RECT  0.165 -0.235 0.465 1.215 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.860 3.685 5.040 4.155 ;
        RECT  4.480 3.250 4.860 4.155 ;
        RECT  3.430 3.685 4.480 4.155 ;
        RECT  3.050 3.250 3.430 4.155 ;
        RECT  1.990 3.685 3.050 4.155 ;
        RECT  1.610 3.250 1.990 4.155 ;
        RECT  0.555 3.685 1.610 4.155 ;
        RECT  0.175 2.630 0.555 4.155 ;
        RECT  0.000 3.685 0.175 4.155 ;
        END
    END VDD
END ND3D2BWP7T

MACRO ND3D3BWP7T
    CLASS CORE ;
    FOREIGN ND3D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 4.6368 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.715 2.380 6.945 3.440 ;
        RECT  5.505 2.380 6.715 2.730 ;
        RECT  5.275 2.380 5.505 3.440 ;
        RECT  4.065 2.380 5.275 2.730 ;
        RECT  3.835 2.380 4.065 3.440 ;
        RECT  2.625 2.380 3.835 2.730 ;
        RECT  2.400 2.380 2.625 3.440 ;
        RECT  2.395 1.020 2.400 3.440 ;
        RECT  1.560 1.020 2.395 2.730 ;
        RECT  0.530 1.020 1.560 1.370 ;
        RECT  1.185 2.390 1.560 2.730 ;
        RECT  0.955 2.390 1.185 3.440 ;
        RECT  0.170 0.490 0.530 1.370 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 1.715 6.480 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.860 1.715 4.320 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.715 1.155 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.015 -0.235 7.280 0.235 ;
        RECT  6.635 -0.235 7.015 1.195 ;
        RECT  5.560 -0.235 6.635 0.235 ;
        RECT  5.215 -0.235 5.560 0.775 ;
        RECT  0.000 -0.235 5.215 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.295 3.685 7.280 4.155 ;
        RECT  5.915 2.960 6.295 4.155 ;
        RECT  4.865 3.685 5.915 4.155 ;
        RECT  4.485 2.960 4.865 4.155 ;
        RECT  3.425 3.685 4.485 4.155 ;
        RECT  3.045 2.960 3.425 4.155 ;
        RECT  1.985 3.685 3.045 4.155 ;
        RECT  1.605 2.960 1.985 4.155 ;
        RECT  0.545 3.685 1.605 4.155 ;
        RECT  0.165 2.535 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.940 0.495 6.280 1.250 ;
        RECT  4.840 1.005 5.940 1.250 ;
        RECT  4.495 0.495 4.840 1.250 ;
        RECT  3.060 1.020 4.495 1.250 ;
        RECT  0.900 0.495 4.120 0.725 ;
    END
END ND3D3BWP7T

MACRO ND3D4BWP7T
    CLASS CORE ;
    FOREIGN ND3D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.5188 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.160 2.380 8.390 3.240 ;
        RECT  6.950 2.380 8.160 2.730 ;
        RECT  6.720 2.380 6.950 3.240 ;
        RECT  5.510 2.380 6.720 2.730 ;
        RECT  5.280 2.380 5.510 3.240 ;
        RECT  4.070 2.380 5.280 2.730 ;
        RECT  3.840 2.380 4.070 3.240 ;
        RECT  2.970 2.380 3.840 2.730 ;
        RECT  2.630 1.015 2.970 2.730 ;
        RECT  2.400 1.015 2.630 3.240 ;
        RECT  2.070 1.015 2.400 2.730 ;
        RECT  0.905 1.015 2.070 1.365 ;
        RECT  1.190 2.380 2.070 2.730 ;
        RECT  0.960 2.380 1.190 3.240 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.545 1.715 9.125 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.675 1.715 5.695 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.715 1.770 1.945 ;
        RECT  0.140 1.715 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.205 -0.235 10.080 0.235 ;
        RECT  8.805 -0.235 9.205 0.730 ;
        RECT  7.765 -0.235 8.805 0.235 ;
        RECT  7.365 -0.235 7.765 0.730 ;
        RECT  0.000 -0.235 7.365 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.180 3.685 10.080 4.155 ;
        RECT  8.800 2.510 9.180 4.155 ;
        RECT  7.740 3.685 8.800 4.155 ;
        RECT  7.360 2.960 7.740 4.155 ;
        RECT  6.310 3.685 7.360 4.155 ;
        RECT  5.930 2.960 6.310 4.155 ;
        RECT  4.870 3.685 5.930 4.155 ;
        RECT  4.490 2.960 4.870 4.155 ;
        RECT  3.430 3.685 4.490 4.155 ;
        RECT  3.050 2.960 3.430 4.155 ;
        RECT  1.990 3.685 3.050 4.155 ;
        RECT  1.610 2.960 1.990 4.155 ;
        RECT  0.520 3.685 1.610 4.155 ;
        RECT  0.180 2.525 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.160 2.380 8.390 3.240 ;
        RECT  6.950 2.380 8.160 2.730 ;
        RECT  6.720 2.380 6.950 3.240 ;
        RECT  5.510 2.380 6.720 2.730 ;
        RECT  5.280 2.380 5.510 3.240 ;
        RECT  4.070 2.380 5.280 2.730 ;
        RECT  3.840 2.380 4.070 3.240 ;
        RECT  3.170 2.380 3.840 2.730 ;
        RECT  0.905 1.015 1.870 1.365 ;
        RECT  1.190 2.380 1.870 2.730 ;
        RECT  0.960 2.380 1.190 3.240 ;
        RECT  9.560 0.495 9.900 1.250 ;
        RECT  8.460 1.005 9.560 1.250 ;
        RECT  8.120 0.495 8.460 1.250 ;
        RECT  3.785 1.020 8.120 1.250 ;
        RECT  0.470 0.465 6.295 0.725 ;
        RECT  0.240 0.465 0.470 1.305 ;
    END
END ND3D4BWP7T

MACRO ND4D0BWP7T
    CLASS CORE ;
    FOREIGN ND4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.0101 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.485 3.220 2.745 ;
        RECT  2.800 0.485 2.940 0.715 ;
        RECT  0.855 2.515 2.940 2.745 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.675 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.810 0.510 2.100 1.590 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.710 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 -0.235 3.360 0.235 ;
        RECT  0.155 -0.235 0.535 0.715 ;
        RECT  0.000 -0.235 0.155 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.190 3.685 3.360 4.155 ;
        RECT  2.820 3.440 3.190 4.155 ;
        RECT  1.965 3.685 2.820 4.155 ;
        RECT  1.600 3.440 1.965 4.155 ;
        RECT  0.595 3.685 1.600 4.155 ;
        RECT  0.240 3.440 0.595 4.155 ;
        RECT  0.000 3.685 0.240 4.155 ;
        END
    END VDD
END ND4D0BWP7T

MACRO ND4D1BWP7T
    CLASS CORE ;
    FOREIGN ND4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.9596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.010 3.780 2.730 ;
        RECT  3.210 1.010 3.500 1.240 ;
        RECT  2.665 2.450 3.500 2.730 ;
        RECT  2.860 0.530 3.210 1.240 ;
        RECT  2.435 2.450 2.665 3.330 ;
        RECT  1.225 2.450 2.435 2.730 ;
        RECT  0.995 2.450 1.225 3.330 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.210 1.540 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.135 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.675 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.560 -0.235 3.920 0.235 ;
        RECT  0.220 -0.235 0.560 1.215 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 3.685 3.920 4.155 ;
        RECT  3.100 2.960 3.440 4.155 ;
        RECT  2.000 3.685 3.100 4.155 ;
        RECT  1.660 2.960 2.000 4.155 ;
        RECT  0.560 3.685 1.660 4.155 ;
        RECT  0.220 2.505 0.560 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
END ND4D1BWP7T

MACRO ND4D2BWP7T
    CLASS CORE ;
    FOREIGN ND4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.4992 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 2.470 6.210 3.390 ;
        RECT  4.550 2.470 5.980 2.750 ;
        RECT  4.320 2.470 4.550 3.390 ;
        RECT  2.910 2.470 4.320 2.750 ;
        RECT  2.680 2.470 2.910 3.390 ;
        RECT  1.850 2.470 2.680 2.750 ;
        RECT  1.285 1.555 1.850 2.750 ;
        RECT  1.230 0.965 1.285 2.750 ;
        RECT  0.955 0.965 1.230 3.430 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.705 1.715 6.580 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.715 5.025 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.345 1.715 3.220 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.715 0.725 1.945 ;
        RECT  0.140 1.715 0.420 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.235 7.280 0.235 ;
        RECT  5.975 -0.235 6.435 0.795 ;
        RECT  0.000 -0.235 5.975 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.005 3.685 7.280 4.155 ;
        RECT  6.620 2.540 7.005 4.155 ;
        RECT  5.475 3.685 6.620 4.155 ;
        RECT  5.090 2.980 5.475 4.155 ;
        RECT  3.805 3.685 5.090 4.155 ;
        RECT  3.420 2.980 3.805 4.155 ;
        RECT  2.175 3.685 3.420 4.155 ;
        RECT  1.790 2.980 2.175 4.155 ;
        RECT  0.610 3.685 1.790 4.155 ;
        RECT  0.225 3.025 0.610 4.155 ;
        RECT  0.000 3.685 0.225 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.745 0.510 7.085 1.275 ;
        RECT  5.590 1.035 6.745 1.275 ;
        RECT  5.360 0.465 5.590 1.275 ;
        RECT  3.865 0.465 5.360 0.700 ;
        RECT  2.385 0.940 4.925 1.170 ;
        RECT  0.510 0.465 3.445 0.700 ;
        RECT  0.280 0.465 0.510 1.275 ;
    END
END ND4D2BWP7T

MACRO ND4D3BWP7T
    CLASS CORE ;
    FOREIGN ND4D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 6.1409 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.920 2.380 9.150 3.390 ;
        RECT  7.710 2.380 8.920 2.730 ;
        RECT  7.480 2.380 7.710 3.390 ;
        RECT  6.270 2.380 7.480 2.730 ;
        RECT  6.040 2.380 6.270 3.390 ;
        RECT  4.830 2.380 6.040 2.730 ;
        RECT  4.600 2.380 4.830 3.390 ;
        RECT  3.390 2.380 4.600 2.730 ;
        RECT  3.160 2.380 3.390 3.390 ;
        RECT  2.410 2.380 3.160 2.730 ;
        RECT  1.950 0.965 2.410 2.730 ;
        RECT  1.720 0.965 1.950 3.390 ;
        RECT  1.510 0.965 1.720 2.730 ;
        RECT  0.505 0.965 1.510 1.315 ;
        RECT  0.505 2.410 1.510 2.730 ;
        RECT  0.275 0.495 0.505 1.315 ;
        RECT  0.275 2.410 0.505 3.390 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.265 1.715 8.645 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.105 1.715 6.485 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.715 4.265 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.715 1.280 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.240 -0.235 9.520 0.235 ;
        RECT  8.860 -0.235 9.240 1.175 ;
        RECT  7.790 -0.235 8.860 0.235 ;
        RECT  7.410 -0.235 7.790 0.785 ;
        RECT  0.000 -0.235 7.410 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.500 3.685 9.520 4.155 ;
        RECT  8.120 2.960 8.500 4.155 ;
        RECT  7.060 3.685 8.120 4.155 ;
        RECT  6.680 2.960 7.060 4.155 ;
        RECT  5.620 3.685 6.680 4.155 ;
        RECT  5.240 2.960 5.620 4.155 ;
        RECT  4.180 3.685 5.240 4.155 ;
        RECT  3.800 2.960 4.180 4.155 ;
        RECT  2.740 3.685 3.800 4.155 ;
        RECT  2.360 2.960 2.740 4.155 ;
        RECT  1.300 3.685 2.360 4.155 ;
        RECT  0.920 2.960 1.300 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.920 2.380 9.150 3.390 ;
        RECT  7.710 2.380 8.920 2.730 ;
        RECT  7.480 2.380 7.710 3.390 ;
        RECT  6.270 2.380 7.480 2.730 ;
        RECT  6.040 2.380 6.270 3.390 ;
        RECT  4.830 2.380 6.040 2.730 ;
        RECT  4.600 2.380 4.830 3.390 ;
        RECT  3.390 2.380 4.600 2.730 ;
        RECT  3.160 2.380 3.390 3.390 ;
        RECT  2.610 2.380 3.160 2.730 ;
        RECT  0.505 0.965 1.310 1.315 ;
        RECT  0.505 2.410 1.310 2.730 ;
        RECT  0.275 0.495 0.505 1.315 ;
        RECT  0.275 2.410 0.505 3.390 ;
        RECT  8.200 0.495 8.430 1.320 ;
        RECT  6.990 1.020 8.200 1.320 ;
        RECT  6.760 0.490 6.990 1.320 ;
        RECT  5.185 0.490 6.760 0.720 ;
        RECT  4.830 1.020 6.325 1.250 ;
        RECT  4.600 0.495 4.830 1.250 ;
        RECT  3.105 1.020 4.600 1.250 ;
        RECT  0.945 0.490 4.165 0.720 ;
    END
END ND4D3BWP7T

MACRO ND4D4BWP7T
    CLASS CORE ;
    FOREIGN ND4D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 6.9962 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.695 2.430 11.925 3.390 ;
        RECT  10.485 2.430 11.695 2.780 ;
        RECT  10.255 2.430 10.485 3.390 ;
        RECT  9.045 2.430 10.255 2.780 ;
        RECT  8.815 2.430 9.045 3.390 ;
        RECT  7.605 2.430 8.815 2.780 ;
        RECT  7.375 2.430 7.605 3.390 ;
        RECT  5.505 2.430 7.375 2.780 ;
        RECT  5.275 2.430 5.505 3.390 ;
        RECT  4.065 2.430 5.275 2.780 ;
        RECT  3.835 2.430 4.065 3.390 ;
        RECT  2.970 2.430 3.835 2.780 ;
        RECT  2.625 1.020 2.970 2.780 ;
        RECT  2.395 1.020 2.625 3.390 ;
        RECT  2.070 1.020 2.395 2.780 ;
        RECT  0.895 1.020 2.070 1.370 ;
        RECT  1.185 2.430 2.070 2.780 ;
        RECT  0.955 2.430 1.185 3.390 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.460 1.770 12.740 2.750 ;
        RECT  10.045 1.770 12.460 2.190 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.185 1.770 9.205 2.190 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 1.7046 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.845 1.770 4.900 2.190 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.680 1.580 2.150 ;
        RECT  0.140 1.210 0.420 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.980 -0.235 12.880 0.235 ;
        RECT  11.640 -0.235 11.980 0.785 ;
        RECT  10.540 -0.235 11.640 0.235 ;
        RECT  10.200 -0.235 10.540 0.785 ;
        RECT  0.000 -0.235 10.200 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.700 3.685 12.880 4.155 ;
        RECT  12.360 3.025 12.700 4.155 ;
        RECT  11.260 3.685 12.360 4.155 ;
        RECT  10.920 3.025 11.260 4.155 ;
        RECT  9.820 3.685 10.920 4.155 ;
        RECT  9.480 3.025 9.820 4.155 ;
        RECT  8.380 3.685 9.480 4.155 ;
        RECT  8.040 3.025 8.380 4.155 ;
        RECT  6.940 3.685 8.040 4.155 ;
        RECT  6.600 3.025 6.940 4.155 ;
        RECT  6.280 3.685 6.600 4.155 ;
        RECT  5.940 3.025 6.280 4.155 ;
        RECT  4.840 3.685 5.940 4.155 ;
        RECT  4.500 3.025 4.840 4.155 ;
        RECT  3.400 3.685 4.500 4.155 ;
        RECT  3.060 3.025 3.400 4.155 ;
        RECT  1.960 3.685 3.060 4.155 ;
        RECT  1.620 3.025 1.960 4.155 ;
        RECT  0.520 3.685 1.620 4.155 ;
        RECT  0.180 2.510 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.695 2.430 11.925 3.390 ;
        RECT  10.485 2.430 11.695 2.780 ;
        RECT  10.255 2.430 10.485 3.390 ;
        RECT  9.045 2.430 10.255 2.780 ;
        RECT  8.815 2.430 9.045 3.390 ;
        RECT  7.605 2.430 8.815 2.780 ;
        RECT  7.375 2.430 7.605 3.390 ;
        RECT  5.505 2.430 7.375 2.780 ;
        RECT  5.275 2.430 5.505 3.390 ;
        RECT  4.065 2.430 5.275 2.780 ;
        RECT  3.835 2.430 4.065 3.390 ;
        RECT  3.170 2.430 3.835 2.780 ;
        RECT  0.895 1.020 1.870 1.370 ;
        RECT  1.185 2.430 1.870 2.780 ;
        RECT  0.955 2.430 1.185 3.390 ;
        RECT  12.415 0.695 12.645 1.250 ;
        RECT  11.205 1.020 12.415 1.250 ;
        RECT  10.975 0.495 11.205 1.250 ;
        RECT  9.765 1.020 10.975 1.250 ;
        RECT  9.535 0.465 9.765 1.250 ;
        RECT  6.600 0.465 9.535 0.695 ;
        RECT  6.850 0.925 9.130 1.155 ;
        RECT  6.620 0.925 6.850 1.775 ;
        RECT  5.750 1.545 6.620 1.775 ;
        RECT  5.995 0.550 6.225 1.315 ;
        RECT  0.180 0.550 5.995 0.780 ;
        RECT  5.520 1.020 5.750 1.775 ;
        RECT  3.775 1.020 5.520 1.250 ;
    END
END ND4D4BWP7T

MACRO NR2D0BWP7T
    CLASS CORE ;
    FOREIGN NR2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6399 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 3.255 ;
        RECT  1.225 1.210 1.820 1.490 ;
        RECT  1.540 3.025 1.820 3.255 ;
        RECT  0.995 0.570 1.225 1.490 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.770 1.540 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.040 -0.235 2.240 0.235 ;
        RECT  1.660 -0.235 2.040 0.855 ;
        RECT  0.600 -0.235 1.660 0.235 ;
        RECT  0.220 -0.235 0.600 0.855 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.560 3.685 2.240 4.155 ;
        RECT  0.220 3.025 0.560 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
END NR2D0BWP7T

MACRO NR2D1BWP7T
    CLASS CORE ;
    FOREIGN NR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 2.505 1.880 3.255 ;
        RECT  1.265 1.165 1.540 3.255 ;
        RECT  1.260 0.495 1.265 3.255 ;
        RECT  1.035 0.495 1.260 1.435 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.715 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 1.210 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.040 -0.235 2.240 0.235 ;
        RECT  1.700 -0.235 2.040 0.915 ;
        RECT  0.565 -0.235 1.700 0.235 ;
        RECT  0.210 -0.235 0.565 1.200 ;
        RECT  0.000 -0.235 0.210 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.590 3.685 2.240 4.155 ;
        RECT  0.210 2.495 0.590 4.155 ;
        RECT  0.000 3.685 0.210 4.155 ;
        END
    END VDD
END NR2D1BWP7T

MACRO NR2D1P5BWP7T
    CLASS CORE ;
    FOREIGN NR2D1P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.3662 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.415 0.465 2.645 1.350 ;
        RECT  2.100 1.070 2.415 1.350 ;
        RECT  1.820 1.070 2.100 2.870 ;
        RECT  1.185 1.070 1.820 1.350 ;
        RECT  1.500 2.640 1.820 2.870 ;
        RECT  0.955 0.500 1.185 1.350 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.6408 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 1.600 3.125 1.980 ;
        RECT  2.580 1.740 2.895 1.980 ;
        RECT  2.340 1.740 2.580 3.340 ;
        RECT  1.080 3.100 2.340 3.340 ;
        RECT  0.840 2.660 1.080 3.340 ;
        RECT  0.450 2.660 0.840 2.900 ;
        RECT  0.140 1.210 0.450 2.900 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6408 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.660 1.545 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 -0.235 3.920 0.235 ;
        RECT  3.080 -0.235 3.460 0.710 ;
        RECT  2.000 -0.235 3.080 0.235 ;
        RECT  1.620 -0.235 2.000 0.710 ;
        RECT  0.560 -0.235 1.620 0.235 ;
        RECT  0.180 -0.235 0.560 0.845 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 3.685 3.920 4.155 ;
        RECT  3.060 2.640 3.440 4.155 ;
        RECT  0.560 3.685 3.060 4.155 ;
        RECT  0.180 3.155 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
END NR2D1P5BWP7T

MACRO NR2D2BWP7T
    CLASS CORE ;
    FOREIGN NR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8198 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.885 1.040 3.530 2.345 ;
        RECT  2.805 1.040 2.885 2.745 ;
        RECT  2.630 0.490 2.805 2.745 ;
        RECT  2.575 0.490 2.630 1.320 ;
        RECT  2.520 2.515 2.630 2.745 ;
        RECT  1.225 1.040 2.575 1.320 ;
        RECT  0.995 0.490 1.225 1.320 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.985 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.715 2.400 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.620 -0.235 3.920 0.235 ;
        RECT  3.240 -0.235 3.620 0.810 ;
        RECT  2.110 -0.235 3.240 0.235 ;
        RECT  1.730 -0.235 2.110 0.810 ;
        RECT  0.560 -0.235 1.730 0.235 ;
        RECT  0.220 -0.235 0.560 1.185 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 3.685 3.920 4.155 ;
        RECT  0.940 2.910 1.280 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.240 2.690 3.580 3.400 ;
        RECT  2.025 3.160 3.240 3.400 ;
        RECT  1.795 2.380 2.025 3.400 ;
        RECT  0.505 2.380 1.795 2.620 ;
        RECT  0.275 2.380 0.505 3.335 ;
    END
END NR2D2BWP7T

MACRO NR2D2P5BWP7T
    CLASS CORE ;
    FOREIGN NR2D2P5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5428 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 1.015 4.900 3.395 ;
        RECT  1.560 1.015 4.575 1.255 ;
        RECT  4.485 2.585 4.575 3.395 ;
        RECT  1.560 2.530 1.840 2.760 ;
        RECT  1.320 1.015 1.560 2.760 ;
        RECT  1.185 1.015 1.320 1.275 ;
        RECT  0.955 0.465 1.185 1.275 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.580 2.010 3.540 2.240 ;
        RECT  2.340 2.010 2.580 3.230 ;
        RECT  1.080 2.990 2.340 3.230 ;
        RECT  0.840 1.910 1.080 3.230 ;
        RECT  0.450 1.910 0.840 2.150 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.0656 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.495 4.345 2.150 ;
        RECT  2.100 1.495 4.060 1.725 ;
        RECT  1.820 1.495 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 -0.235 5.040 0.235 ;
        RECT  3.040 -0.235 3.500 0.785 ;
        RECT  2.050 -0.235 3.040 0.235 ;
        RECT  1.590 -0.235 2.050 0.785 ;
        RECT  0.560 -0.235 1.590 0.235 ;
        RECT  0.180 -0.235 0.560 0.895 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 3.685 5.040 4.155 ;
        RECT  2.920 2.710 3.300 4.155 ;
        RECT  0.560 3.685 2.920 4.155 ;
        RECT  0.180 2.580 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
END NR2D2P5BWP7T

MACRO NR2D3BWP7T
    CLASS CORE ;
    FOREIGN NR2D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0174 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 2.465 4.805 3.295 ;
        RECT  4.090 2.465 4.575 2.765 ;
        RECT  3.855 0.495 4.090 2.765 ;
        RECT  3.190 1.040 3.855 2.765 ;
        RECT  2.645 1.040 3.190 1.340 ;
        RECT  3.080 2.465 3.190 2.765 ;
        RECT  2.415 0.495 2.645 1.340 ;
        RECT  1.205 1.040 2.415 1.340 ;
        RECT  0.975 0.495 1.205 1.340 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 1.660 2.100 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.2798 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.210 4.900 2.150 ;
        RECT  4.320 1.660 4.620 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 -0.235 5.040 0.235 ;
        RECT  4.480 -0.235 4.880 0.980 ;
        RECT  3.440 -0.235 4.480 0.235 ;
        RECT  3.060 -0.235 3.440 0.810 ;
        RECT  2.020 -0.235 3.060 0.235 ;
        RECT  1.640 -0.235 2.020 0.810 ;
        RECT  0.580 -0.235 1.640 0.235 ;
        RECT  0.200 -0.235 0.580 1.215 ;
        RECT  0.000 -0.235 0.200 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.020 3.685 5.040 4.155 ;
        RECT  1.640 2.935 2.020 4.155 ;
        RECT  0.580 3.685 1.640 4.155 ;
        RECT  0.200 2.575 0.580 4.155 ;
        RECT  0.000 3.685 0.200 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.645 3.105 4.140 3.335 ;
        RECT  2.415 2.475 2.645 3.335 ;
        RECT  1.205 2.475 2.415 2.705 ;
        RECT  0.975 2.475 1.205 3.335 ;
    END
END NR2D3BWP7T

MACRO NR2D4BWP7T
    CLASS CORE ;
    FOREIGN NR2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.6396 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.650 2.550 5.600 2.780 ;
        RECT  5.315 0.495 5.545 1.360 ;
        RECT  4.650 1.040 5.315 1.360 ;
        RECT  4.105 1.040 4.650 2.780 ;
        RECT  3.875 0.495 4.105 2.780 ;
        RECT  3.750 1.040 3.875 2.780 ;
        RECT  2.665 1.040 3.750 1.360 ;
        RECT  2.435 0.495 2.665 1.360 ;
        RECT  1.225 1.040 2.435 1.360 ;
        RECT  0.995 0.495 1.225 1.360 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.715 2.930 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.7064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.900 1.715 6.020 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.320 -0.235 6.720 0.235 ;
        RECT  5.980 -0.235 6.320 1.190 ;
        RECT  4.900 -0.235 5.980 0.235 ;
        RECT  4.520 -0.235 4.900 0.810 ;
        RECT  3.440 -0.235 4.520 0.235 ;
        RECT  3.100 -0.235 3.440 0.810 ;
        RECT  2.000 -0.235 3.100 0.235 ;
        RECT  1.660 -0.235 2.000 0.810 ;
        RECT  0.560 -0.235 1.660 0.235 ;
        RECT  0.220 -0.235 0.560 1.190 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 3.685 6.720 4.155 ;
        RECT  2.380 2.990 2.760 4.155 ;
        RECT  1.320 3.685 2.380 4.155 ;
        RECT  0.940 2.990 1.320 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.850 2.550 5.600 2.780 ;
        RECT  5.315 0.495 5.545 1.360 ;
        RECT  4.850 1.040 5.315 1.360 ;
        RECT  2.665 1.040 3.550 1.360 ;
        RECT  2.435 0.495 2.665 1.360 ;
        RECT  1.225 1.040 2.435 1.360 ;
        RECT  0.995 0.495 1.225 1.360 ;
        RECT  6.035 2.480 6.265 3.290 ;
        RECT  3.385 3.060 6.035 3.290 ;
        RECT  3.155 2.480 3.385 3.290 ;
        RECT  1.945 2.480 3.155 2.760 ;
        RECT  1.715 2.480 1.945 3.290 ;
        RECT  0.505 2.480 1.715 2.760 ;
        RECT  0.275 2.480 0.505 3.290 ;
    END
END NR2D4BWP7T

MACRO NR2D5BWP7T
    CLASS CORE ;
    FOREIGN NR2D5BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.6690 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.815 0.495 8.045 1.485 ;
        RECT  7.815 2.420 8.045 3.230 ;
        RECT  6.525 1.135 7.815 1.485 ;
        RECT  5.770 2.420 7.815 2.770 ;
        RECT  6.295 0.495 6.525 1.485 ;
        RECT  5.770 1.135 6.295 1.485 ;
        RECT  5.025 1.135 5.770 2.770 ;
        RECT  4.870 0.495 5.025 2.770 ;
        RECT  4.795 0.495 4.870 1.485 ;
        RECT  4.740 2.420 4.870 2.770 ;
        RECT  3.505 1.135 4.795 1.485 ;
        RECT  3.275 0.495 3.505 1.485 ;
        RECT  2.005 1.135 3.275 1.485 ;
        RECT  1.775 0.495 2.005 1.485 ;
        RECT  0.485 1.135 1.775 1.485 ;
        RECT  0.255 0.495 0.485 1.485 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 2.1330 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.715 3.570 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.1330 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.160 1.715 7.440 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.350 -0.235 8.400 0.235 ;
        RECT  7.010 -0.235 7.350 0.905 ;
        RECT  5.830 -0.235 7.010 0.235 ;
        RECT  5.490 -0.235 5.830 0.905 ;
        RECT  4.320 -0.235 5.490 0.235 ;
        RECT  3.980 -0.235 4.320 0.905 ;
        RECT  2.810 -0.235 3.980 0.235 ;
        RECT  2.470 -0.235 2.810 0.905 ;
        RECT  1.350 -0.235 2.470 0.235 ;
        RECT  0.970 -0.235 1.350 0.905 ;
        RECT  0.000 -0.235 0.970 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.560 3.685 8.400 4.155 ;
        RECT  3.220 2.960 3.560 4.155 ;
        RECT  2.060 3.685 3.220 4.155 ;
        RECT  1.680 2.960 2.060 4.155 ;
        RECT  0.495 3.685 1.680 4.155 ;
        RECT  0.240 2.245 0.495 4.155 ;
        RECT  0.000 3.685 0.240 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.815 0.495 8.045 1.485 ;
        RECT  7.815 2.420 8.045 3.230 ;
        RECT  6.525 1.135 7.815 1.485 ;
        RECT  5.970 2.420 7.815 2.770 ;
        RECT  6.295 0.495 6.525 1.485 ;
        RECT  5.970 1.135 6.295 1.485 ;
        RECT  3.505 1.135 4.670 1.485 ;
        RECT  3.275 0.495 3.505 1.485 ;
        RECT  2.005 1.135 3.275 1.485 ;
        RECT  1.775 0.495 2.005 1.485 ;
        RECT  0.485 1.135 1.775 1.485 ;
        RECT  0.255 0.495 0.485 1.485 ;
        RECT  4.265 3.030 7.360 3.260 ;
        RECT  4.035 2.450 4.265 3.260 ;
        RECT  2.745 2.450 4.035 2.730 ;
        RECT  2.515 2.450 2.745 3.320 ;
        RECT  1.225 2.450 2.515 2.730 ;
        RECT  0.995 2.450 1.225 3.320 ;
    END
END NR2D5BWP7T

MACRO NR2D6BWP7T
    CLASS CORE ;
    FOREIGN NR2D6BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.5394 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.330 2.455 8.620 2.805 ;
        RECT  8.195 0.475 8.425 1.440 ;
        RECT  6.985 1.120 8.195 1.440 ;
        RECT  6.755 0.475 6.985 1.440 ;
        RECT  6.330 1.120 6.755 1.440 ;
        RECT  5.545 1.120 6.330 2.805 ;
        RECT  5.430 0.475 5.545 2.805 ;
        RECT  5.315 0.475 5.430 1.440 ;
        RECT  5.260 2.455 5.430 2.805 ;
        RECT  4.105 1.120 5.315 1.440 ;
        RECT  3.875 0.475 4.105 1.440 ;
        RECT  2.665 1.120 3.875 1.440 ;
        RECT  2.435 0.475 2.665 1.440 ;
        RECT  1.225 1.120 2.435 1.440 ;
        RECT  0.995 0.475 1.225 1.440 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 2.5596 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.705 1.715 4.335 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.5596 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.775 1.715 8.525 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.260 -0.235 9.520 0.235 ;
        RECT  8.880 -0.235 9.260 1.230 ;
        RECT  7.800 -0.235 8.880 0.235 ;
        RECT  7.420 -0.235 7.800 0.865 ;
        RECT  6.360 -0.235 7.420 0.235 ;
        RECT  5.980 -0.235 6.360 0.865 ;
        RECT  4.920 -0.235 5.980 0.235 ;
        RECT  4.540 -0.235 4.920 0.865 ;
        RECT  3.480 -0.235 4.540 0.235 ;
        RECT  3.100 -0.235 3.480 0.865 ;
        RECT  2.040 -0.235 3.100 0.235 ;
        RECT  1.660 -0.235 2.040 0.865 ;
        RECT  0.560 -0.235 1.660 0.235 ;
        RECT  0.180 -0.235 0.560 1.205 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 3.685 9.520 4.155 ;
        RECT  3.820 3.000 4.200 4.155 ;
        RECT  2.720 3.685 3.820 4.155 ;
        RECT  2.340 3.000 2.720 4.155 ;
        RECT  1.280 3.685 2.340 4.155 ;
        RECT  0.900 3.000 1.280 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.530 2.455 8.620 2.805 ;
        RECT  8.195 0.475 8.425 1.440 ;
        RECT  6.985 1.120 8.195 1.440 ;
        RECT  6.755 0.475 6.985 1.440 ;
        RECT  6.530 1.120 6.755 1.440 ;
        RECT  4.105 1.120 5.230 1.440 ;
        RECT  3.875 0.475 4.105 1.440 ;
        RECT  2.665 1.120 3.875 1.440 ;
        RECT  2.435 0.475 2.665 1.440 ;
        RECT  1.225 1.120 2.435 1.440 ;
        RECT  0.995 0.475 1.225 1.440 ;
        RECT  8.955 2.470 9.185 3.280 ;
        RECT  4.825 3.045 8.955 3.280 ;
        RECT  4.595 2.460 4.825 3.280 ;
        RECT  3.385 2.460 4.595 2.760 ;
        RECT  3.155 2.460 3.385 3.280 ;
        RECT  1.925 2.460 3.155 2.760 ;
        RECT  1.695 2.460 1.925 3.280 ;
        RECT  0.465 2.460 1.695 2.760 ;
        RECT  0.235 2.460 0.465 3.280 ;
    END
END NR2D6BWP7T

MACRO NR2D8BWP7T
    CLASS CORE ;
    FOREIGN NR2D8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.320 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 7.2792 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.450 2.450 11.365 2.770 ;
        RECT  11.080 0.495 11.310 1.440 ;
        RECT  9.870 1.120 11.080 1.440 ;
        RECT  9.640 0.495 9.870 1.440 ;
        RECT  8.430 1.120 9.640 1.440 ;
        RECT  8.200 0.495 8.430 1.440 ;
        RECT  7.450 1.120 8.200 1.440 ;
        RECT  6.990 1.120 7.450 2.770 ;
        RECT  6.760 0.495 6.990 2.770 ;
        RECT  6.550 1.120 6.760 2.770 ;
        RECT  5.550 1.120 6.550 1.440 ;
        RECT  5.320 0.495 5.550 1.440 ;
        RECT  4.110 1.120 5.320 1.440 ;
        RECT  3.880 0.495 4.110 1.440 ;
        RECT  2.670 1.120 3.880 1.440 ;
        RECT  2.440 0.495 2.670 1.440 ;
        RECT  1.230 1.120 2.440 1.440 ;
        RECT  1.000 0.495 1.230 1.440 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 3.4128 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.755 1.715 5.795 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 3.4128 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.950 1.715 11.635 2.110 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.105 -0.235 12.320 0.235 ;
        RECT  11.700 -0.235 12.105 1.185 ;
        RECT  10.685 -0.235 11.700 0.235 ;
        RECT  10.300 -0.235 10.685 0.865 ;
        RECT  9.245 -0.235 10.300 0.235 ;
        RECT  8.860 -0.235 9.245 0.865 ;
        RECT  7.805 -0.235 8.860 0.235 ;
        RECT  7.420 -0.235 7.805 0.865 ;
        RECT  6.365 -0.235 7.420 0.235 ;
        RECT  5.980 -0.235 6.365 0.865 ;
        RECT  4.925 -0.235 5.980 0.235 ;
        RECT  4.540 -0.235 4.925 0.865 ;
        RECT  3.445 -0.235 4.540 0.235 ;
        RECT  3.100 -0.235 3.445 0.865 ;
        RECT  2.005 -0.235 3.100 0.235 ;
        RECT  1.660 -0.235 2.005 0.865 ;
        RECT  0.575 -0.235 1.660 0.235 ;
        RECT  0.215 -0.235 0.575 1.185 ;
        RECT  0.000 -0.235 0.215 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.640 3.685 12.320 4.155 ;
        RECT  5.260 3.155 5.640 4.155 ;
        RECT  4.200 3.685 5.260 4.155 ;
        RECT  3.820 3.155 4.200 4.155 ;
        RECT  2.760 3.685 3.820 4.155 ;
        RECT  2.380 3.155 2.760 4.155 ;
        RECT  1.320 3.685 2.380 4.155 ;
        RECT  0.940 3.155 1.320 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.650 2.450 11.365 2.770 ;
        RECT  11.080 0.495 11.310 1.440 ;
        RECT  9.870 1.120 11.080 1.440 ;
        RECT  9.640 0.495 9.870 1.440 ;
        RECT  8.430 1.120 9.640 1.440 ;
        RECT  8.200 0.495 8.430 1.440 ;
        RECT  7.650 1.120 8.200 1.440 ;
        RECT  5.550 1.120 6.350 1.440 ;
        RECT  5.320 0.495 5.550 1.440 ;
        RECT  4.110 1.120 5.320 1.440 ;
        RECT  3.880 0.495 4.110 1.440 ;
        RECT  2.670 1.120 3.880 1.440 ;
        RECT  2.440 0.495 2.670 1.440 ;
        RECT  1.230 1.120 2.440 1.440 ;
        RECT  1.000 0.495 1.230 1.440 ;
        RECT  11.800 2.505 12.030 3.315 ;
        RECT  6.270 3.085 11.800 3.315 ;
        RECT  6.040 2.470 6.270 3.315 ;
        RECT  4.830 2.470 6.040 2.770 ;
        RECT  4.600 2.470 4.830 3.280 ;
        RECT  3.390 2.470 4.600 2.770 ;
        RECT  3.160 2.470 3.390 3.280 ;
        RECT  1.950 2.470 3.160 2.770 ;
        RECT  1.720 2.470 1.950 3.280 ;
        RECT  0.510 2.470 1.720 2.770 ;
        RECT  0.280 2.470 0.510 3.280 ;
    END
END NR2D8BWP7T

MACRO NR2XD0BWP7T
    CLASS CORE ;
    FOREIGN NR2XD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.0098 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.095 2.100 3.310 ;
        RECT  1.290 1.095 1.820 1.335 ;
        RECT  1.655 2.500 1.820 3.310 ;
        RECT  1.050 0.480 1.290 1.335 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.735 1.560 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 -0.235 2.240 0.235 ;
        RECT  1.720 -0.235 2.100 0.725 ;
        RECT  0.660 -0.235 1.720 0.235 ;
        RECT  0.280 -0.235 0.660 0.745 ;
        RECT  0.000 -0.235 0.280 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.660 3.685 2.240 4.155 ;
        RECT  0.280 2.545 0.660 4.155 ;
        RECT  0.000 3.685 0.280 4.155 ;
        END
    END VDD
END NR2XD0BWP7T

MACRO NR2XD1BWP7T
    CLASS CORE ;
    FOREIGN NR2XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.655 2.245 2.885 2.975 ;
        RECT  2.100 2.245 2.655 2.475 ;
        RECT  2.100 0.495 2.165 1.400 ;
        RECT  1.935 0.495 2.100 2.475 ;
        RECT  1.820 1.170 1.935 2.475 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.680 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        RECT  2.700 1.680 3.500 1.910 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.960 -0.235 3.920 0.235 ;
        RECT  2.580 -0.235 2.960 1.200 ;
        RECT  1.450 -0.235 2.580 0.235 ;
        RECT  1.210 -0.235 1.450 1.255 ;
        RECT  0.000 -0.235 1.210 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.530 3.685 3.920 4.155 ;
        RECT  1.150 3.165 1.530 4.155 ;
        RECT  0.000 3.685 1.150 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.375 2.410 3.605 3.455 ;
        RECT  2.220 3.215 3.375 3.455 ;
        RECT  1.880 2.705 2.220 3.455 ;
        RECT  0.725 2.705 1.880 2.935 ;
        RECT  0.495 2.450 0.725 3.415 ;
    END
END NR2XD1BWP7T

MACRO NR2XD2BWP7T
    CLASS CORE ;
    FOREIGN NR2XD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.305 2.225 5.555 2.955 ;
        RECT  4.340 2.225 5.305 2.505 ;
        RECT  4.110 1.075 4.340 2.505 ;
        RECT  4.105 1.075 4.110 2.955 ;
        RECT  4.060 0.495 4.105 2.955 ;
        RECT  3.875 0.495 4.060 1.355 ;
        RECT  3.865 2.225 4.060 2.955 ;
        RECT  2.665 1.075 3.875 1.355 ;
        RECT  2.435 0.495 2.665 1.355 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.660 2.930 1.890 ;
        RECT  0.700 0.650 0.980 1.890 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 0.650 6.030 1.945 ;
        RECT  4.615 1.605 5.740 1.945 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.920 -0.235 6.720 0.235 ;
        RECT  4.580 -0.235 4.920 1.240 ;
        RECT  3.460 -0.235 4.580 0.235 ;
        RECT  3.080 -0.235 3.460 0.805 ;
        RECT  2.000 -0.235 3.080 0.235 ;
        RECT  1.660 -0.235 2.000 1.240 ;
        RECT  0.000 -0.235 1.660 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.760 3.685 6.720 4.155 ;
        RECT  2.380 2.875 2.760 4.155 ;
        RECT  1.300 3.685 2.380 4.155 ;
        RECT  0.920 2.875 1.300 4.155 ;
        RECT  0.000 3.685 0.920 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.035 2.420 6.265 3.455 ;
        RECT  4.880 3.225 6.035 3.455 ;
        RECT  4.540 2.735 4.880 3.455 ;
        RECT  3.385 3.225 4.540 3.455 ;
        RECT  3.155 2.250 3.385 3.455 ;
        RECT  1.945 2.250 3.155 2.530 ;
        RECT  1.715 2.250 1.945 3.405 ;
        RECT  0.505 2.250 1.715 2.530 ;
        RECT  0.275 2.250 0.505 3.405 ;
    END
END NR2XD2BWP7T

MACRO NR2XD3BWP7T
    CLASS CORE ;
    FOREIGN NR2XD3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 4.3308 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.635 0.485 7.865 1.245 ;
        RECT  7.635 2.380 7.865 3.425 ;
        RECT  6.425 0.945 7.635 1.245 ;
        RECT  5.770 2.380 7.635 2.680 ;
        RECT  6.195 0.485 6.425 1.245 ;
        RECT  5.770 0.945 6.195 1.245 ;
        RECT  4.985 0.945 5.770 2.680 ;
        RECT  4.870 0.485 4.985 2.680 ;
        RECT  4.755 0.485 4.870 1.245 ;
        RECT  4.700 2.380 4.870 2.680 ;
        RECT  3.545 0.945 4.755 1.245 ;
        RECT  3.315 0.485 3.545 1.245 ;
        RECT  2.105 0.945 3.315 1.245 ;
        RECT  1.875 0.485 2.105 1.245 ;
        RECT  0.665 0.945 1.875 1.245 ;
        RECT  0.435 0.485 0.665 1.245 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 2.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.770 7.700 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.240 -0.235 8.400 0.235 ;
        RECT  6.860 -0.235 7.240 0.710 ;
        RECT  5.780 -0.235 6.860 0.235 ;
        RECT  5.400 -0.235 5.780 0.710 ;
        RECT  4.340 -0.235 5.400 0.235 ;
        RECT  3.960 -0.235 4.340 0.710 ;
        RECT  2.920 -0.235 3.960 0.235 ;
        RECT  2.540 -0.235 2.920 0.710 ;
        RECT  1.470 -0.235 2.540 0.235 ;
        RECT  1.090 -0.235 1.470 0.710 ;
        RECT  0.000 -0.235 1.090 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.600 3.685 8.400 4.155 ;
        RECT  3.260 2.590 3.600 4.155 ;
        RECT  2.160 3.685 3.260 4.155 ;
        RECT  1.820 2.910 2.160 4.155 ;
        RECT  0.660 3.685 1.820 4.155 ;
        RECT  0.280 2.690 0.660 4.155 ;
        RECT  0.000 3.685 0.280 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.265 2.910 7.200 3.140 ;
        RECT  4.035 2.050 4.265 3.345 ;
        RECT  2.825 2.050 4.035 2.330 ;
        RECT  2.595 2.050 2.825 3.330 ;
        RECT  1.385 2.400 2.595 2.680 ;
        RECT  1.155 2.400 1.385 3.340 ;
    END
END NR2XD3BWP7T

MACRO NR2XD4BWP7T
    CLASS CORE ;
    FOREIGN NR2XD4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.200 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.7270 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.445 0.495 10.675 1.305 ;
        RECT  10.445 2.380 10.675 3.240 ;
        RECT  9.235 0.955 10.445 1.305 ;
        RECT  6.890 2.380 10.445 2.730 ;
        RECT  9.005 0.485 9.235 1.305 ;
        RECT  7.795 0.955 9.005 1.305 ;
        RECT  7.565 0.495 7.795 1.305 ;
        RECT  6.890 0.955 7.565 1.305 ;
        RECT  6.355 0.955 6.890 2.730 ;
        RECT  6.125 0.485 6.355 2.730 ;
        RECT  5.990 0.955 6.125 2.730 ;
        RECT  4.915 0.955 5.990 1.305 ;
        RECT  4.685 0.485 4.915 1.305 ;
        RECT  3.475 0.955 4.685 1.305 ;
        RECT  3.245 0.485 3.475 1.305 ;
        RECT  2.035 0.955 3.245 1.305 ;
        RECT  1.805 0.485 2.035 1.305 ;
        RECT  0.595 0.955 1.805 1.305 ;
        RECT  0.365 0.485 0.595 1.305 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 2.6910 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.540 5.065 1.770 ;
        RECT  0.700 1.540 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.6910 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.540 10.500 2.150 ;
        RECT  7.560 1.540 9.660 1.770 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.030 -0.235 11.200 0.235 ;
        RECT  9.650 -0.235 10.030 0.720 ;
        RECT  8.590 -0.235 9.650 0.235 ;
        RECT  8.210 -0.235 8.590 0.720 ;
        RECT  7.150 -0.235 8.210 0.235 ;
        RECT  6.770 -0.235 7.150 0.720 ;
        RECT  5.730 -0.235 6.770 0.235 ;
        RECT  5.350 -0.235 5.730 0.720 ;
        RECT  4.280 -0.235 5.350 0.235 ;
        RECT  3.900 -0.235 4.280 0.720 ;
        RECT  2.850 -0.235 3.900 0.235 ;
        RECT  2.470 -0.235 2.850 0.720 ;
        RECT  1.400 -0.235 2.470 0.235 ;
        RECT  1.020 -0.235 1.400 0.720 ;
        RECT  0.000 -0.235 1.020 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.970 3.685 11.200 4.155 ;
        RECT  4.630 3.005 4.970 4.155 ;
        RECT  3.550 3.685 4.630 4.155 ;
        RECT  3.170 3.005 3.550 4.155 ;
        RECT  2.090 3.685 3.170 4.155 ;
        RECT  1.750 3.005 2.090 4.155 ;
        RECT  0.670 3.685 1.750 4.155 ;
        RECT  0.290 2.455 0.670 4.155 ;
        RECT  0.000 3.685 0.290 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.445 0.495 10.675 1.305 ;
        RECT  10.445 2.380 10.675 3.240 ;
        RECT  9.235 0.955 10.445 1.305 ;
        RECT  7.090 2.380 10.445 2.730 ;
        RECT  9.005 0.485 9.235 1.305 ;
        RECT  7.795 0.955 9.005 1.305 ;
        RECT  7.565 0.495 7.795 1.305 ;
        RECT  7.090 0.955 7.565 1.305 ;
        RECT  4.915 0.955 5.790 1.305 ;
        RECT  4.685 0.485 4.915 1.305 ;
        RECT  3.475 0.955 4.685 1.305 ;
        RECT  3.245 0.485 3.475 1.305 ;
        RECT  2.035 0.955 3.245 1.305 ;
        RECT  1.805 0.485 2.035 1.305 ;
        RECT  0.595 0.955 1.805 1.305 ;
        RECT  0.365 0.485 0.595 1.305 ;
        RECT  5.635 3.070 10.010 3.350 ;
        RECT  5.405 2.450 5.635 3.350 ;
        RECT  4.195 2.450 5.405 2.730 ;
        RECT  3.965 2.450 4.195 3.320 ;
        RECT  2.755 2.450 3.965 2.730 ;
        RECT  2.525 2.450 2.755 3.320 ;
        RECT  1.315 2.450 2.525 2.730 ;
        RECT  1.085 2.450 1.315 3.320 ;
    END
END NR2XD4BWP7T

MACRO NR2XD8BWP7T
    CLASS CORE ;
    FOREIGN NR2XD8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 10.7424 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.090 0.525 19.320 1.310 ;
        RECT  19.090 2.430 19.320 3.340 ;
        RECT  17.880 0.960 19.090 1.310 ;
        RECT  11.370 2.430 19.090 2.780 ;
        RECT  17.650 0.525 17.880 1.310 ;
        RECT  16.440 0.960 17.650 1.310 ;
        RECT  16.210 0.525 16.440 1.310 ;
        RECT  15.000 0.960 16.210 1.310 ;
        RECT  14.770 0.525 15.000 1.310 ;
        RECT  13.560 0.960 14.770 1.310 ;
        RECT  13.330 0.525 13.560 1.310 ;
        RECT  12.120 0.960 13.330 1.310 ;
        RECT  11.890 0.525 12.120 1.310 ;
        RECT  11.370 0.960 11.890 1.310 ;
        RECT  10.675 0.960 11.370 2.780 ;
        RECT  10.470 0.525 10.675 2.780 ;
        RECT  10.445 0.525 10.470 1.310 ;
        RECT  10.390 2.430 10.470 2.780 ;
        RECT  9.235 0.960 10.445 1.310 ;
        RECT  9.005 0.525 9.235 1.310 ;
        RECT  7.795 0.960 9.005 1.310 ;
        RECT  7.565 0.525 7.795 1.310 ;
        RECT  6.355 0.960 7.565 1.310 ;
        RECT  6.125 0.525 6.355 1.310 ;
        RECT  4.915 0.960 6.125 1.310 ;
        RECT  4.685 0.525 4.915 1.310 ;
        RECT  3.475 0.960 4.685 1.310 ;
        RECT  3.245 0.525 3.475 1.310 ;
        RECT  2.035 0.960 3.245 1.310 ;
        RECT  1.805 0.525 2.035 1.310 ;
        RECT  0.595 0.960 1.805 1.310 ;
        RECT  0.365 0.525 0.595 1.310 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 5.3856 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 1.005 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 5.3856 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.620 1.770 19.460 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.680 -0.235 19.600 0.235 ;
        RECT  18.300 -0.235 18.680 0.730 ;
        RECT  17.250 -0.235 18.300 0.235 ;
        RECT  16.870 -0.235 17.250 0.730 ;
        RECT  15.790 -0.235 16.870 0.235 ;
        RECT  15.410 -0.235 15.790 0.730 ;
        RECT  14.350 -0.235 15.410 0.235 ;
        RECT  13.970 -0.235 14.350 0.730 ;
        RECT  12.910 -0.235 13.970 0.235 ;
        RECT  12.530 -0.235 12.910 0.730 ;
        RECT  11.490 -0.235 12.530 0.235 ;
        RECT  11.110 -0.235 11.490 0.730 ;
        RECT  10.040 -0.235 11.110 0.235 ;
        RECT  9.660 -0.235 10.040 0.730 ;
        RECT  8.590 -0.235 9.660 0.235 ;
        RECT  8.210 -0.235 8.590 0.730 ;
        RECT  7.160 -0.235 8.210 0.235 ;
        RECT  6.780 -0.235 7.160 0.730 ;
        RECT  5.730 -0.235 6.780 0.235 ;
        RECT  5.350 -0.235 5.730 0.730 ;
        RECT  4.280 -0.235 5.350 0.235 ;
        RECT  3.900 -0.235 4.280 0.730 ;
        RECT  2.830 -0.235 3.900 0.235 ;
        RECT  2.450 -0.235 2.830 0.730 ;
        RECT  1.400 -0.235 2.450 0.235 ;
        RECT  1.020 -0.235 1.400 0.730 ;
        RECT  0.000 -0.235 1.020 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.330 3.685 19.600 4.155 ;
        RECT  8.950 2.620 9.330 4.155 ;
        RECT  7.870 3.685 8.950 4.155 ;
        RECT  7.490 2.620 7.870 4.155 ;
        RECT  6.450 3.685 7.490 4.155 ;
        RECT  6.070 2.620 6.450 4.155 ;
        RECT  4.990 3.685 6.070 4.155 ;
        RECT  4.610 2.620 4.990 4.155 ;
        RECT  3.570 3.685 4.610 4.155 ;
        RECT  3.190 2.620 3.570 4.155 ;
        RECT  2.110 3.685 3.190 4.155 ;
        RECT  1.730 2.975 2.110 4.155 ;
        RECT  0.610 3.685 1.730 4.155 ;
        RECT  0.230 2.585 0.610 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.090 0.525 19.320 1.310 ;
        RECT  19.090 2.430 19.320 3.340 ;
        RECT  17.880 0.960 19.090 1.310 ;
        RECT  11.570 2.430 19.090 2.780 ;
        RECT  17.650 0.525 17.880 1.310 ;
        RECT  16.440 0.960 17.650 1.310 ;
        RECT  16.210 0.525 16.440 1.310 ;
        RECT  15.000 0.960 16.210 1.310 ;
        RECT  14.770 0.525 15.000 1.310 ;
        RECT  13.560 0.960 14.770 1.310 ;
        RECT  13.330 0.525 13.560 1.310 ;
        RECT  12.120 0.960 13.330 1.310 ;
        RECT  11.890 0.525 12.120 1.310 ;
        RECT  11.570 0.960 11.890 1.310 ;
        RECT  9.235 0.960 10.270 1.310 ;
        RECT  9.005 0.525 9.235 1.310 ;
        RECT  7.795 0.960 9.005 1.310 ;
        RECT  7.565 0.525 7.795 1.310 ;
        RECT  6.355 0.960 7.565 1.310 ;
        RECT  6.125 0.525 6.355 1.310 ;
        RECT  4.915 0.960 6.125 1.310 ;
        RECT  4.685 0.525 4.915 1.310 ;
        RECT  3.475 0.960 4.685 1.310 ;
        RECT  3.245 0.525 3.475 1.310 ;
        RECT  2.035 0.960 3.245 1.310 ;
        RECT  1.805 0.525 2.035 1.310 ;
        RECT  0.595 0.960 1.805 1.310 ;
        RECT  0.365 0.525 0.595 1.310 ;
        RECT  9.955 3.120 18.755 3.400 ;
        RECT  9.725 2.080 9.955 3.400 ;
        RECT  8.515 2.080 9.725 2.340 ;
        RECT  8.285 2.080 8.515 3.360 ;
        RECT  7.075 2.080 8.285 2.340 ;
        RECT  6.845 2.080 7.075 3.360 ;
        RECT  5.635 2.080 6.845 2.340 ;
        RECT  5.405 2.080 5.635 3.360 ;
        RECT  4.195 2.080 5.405 2.340 ;
        RECT  3.965 2.080 4.195 3.360 ;
        RECT  2.755 2.080 3.965 2.340 ;
        RECT  2.525 2.080 2.755 3.360 ;
        RECT  1.315 2.440 2.525 2.700 ;
        RECT  1.085 2.440 1.315 3.350 ;
    END
END NR2XD8BWP7T

MACRO NR3D0BWP7T
    CLASS CORE ;
    FOREIGN NR3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1676 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.905 2.660 3.170 ;
        RECT  0.900 0.905 2.380 1.135 ;
        RECT  2.105 2.940 2.380 3.170 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.735 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.690 2.100 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.525 -0.235 2.800 0.235 ;
        RECT  0.185 -0.235 0.525 1.135 ;
        RECT  0.000 -0.235 0.185 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 3.685 2.800 4.155 ;
        RECT  0.170 3.025 0.550 4.155 ;
        RECT  0.000 3.685 0.170 4.155 ;
        END
    END VDD
END NR3D0BWP7T

MACRO NR3D1BWP7T
    CLASS CORE ;
    FOREIGN NR3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.7598 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.625 4.340 2.455 ;
        RECT  2.820 0.625 4.060 0.865 ;
        RECT  3.680 2.215 4.060 2.455 ;
        RECT  3.450 2.215 3.680 3.220 ;
        RECT  2.100 2.940 3.450 3.220 ;
        RECT  2.380 0.625 2.820 0.925 ;
        RECT  1.205 0.695 2.380 0.925 ;
        RECT  0.975 0.520 1.205 0.925 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 1.095 3.820 1.490 ;
        RECT  0.980 1.210 3.450 1.490 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.460 1.660 0.700 2.000 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.770 3.360 2.000 ;
        RECT  2.940 1.770 3.220 2.660 ;
        RECT  1.540 2.380 2.940 2.660 ;
        RECT  1.215 1.720 1.540 2.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.770 2.670 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.050 -0.235 4.480 0.235 ;
        RECT  1.670 -0.235 2.050 0.465 ;
        RECT  0.560 -0.235 1.670 0.235 ;
        RECT  0.180 -0.235 0.560 0.985 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.290 3.685 4.480 4.155 ;
        RECT  3.910 2.685 4.290 4.155 ;
        RECT  0.560 3.685 3.910 4.155 ;
        RECT  0.180 2.660 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
END NR3D1BWP7T

MACRO NR3D2BWP7T
    CLASS CORE ;
    FOREIGN NR3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.6750 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.595 2.595 9.825 3.405 ;
        RECT  8.010 2.595 9.595 2.825 ;
        RECT  8.875 0.465 9.105 1.185 ;
        RECT  8.010 0.905 8.875 1.185 ;
        RECT  7.665 0.905 8.010 2.825 ;
        RECT  7.435 0.465 7.665 2.825 ;
        RECT  7.110 0.905 7.435 2.825 ;
        RECT  5.505 0.905 7.110 1.185 ;
        RECT  6.660 2.595 7.110 2.825 ;
        RECT  5.275 0.465 5.505 1.185 ;
        RECT  4.065 0.905 5.275 1.185 ;
        RECT  3.835 0.465 4.065 1.185 ;
        RECT  2.625 0.905 3.835 1.185 ;
        RECT  2.395 0.465 2.625 1.185 ;
        RECT  1.185 0.905 2.395 1.185 ;
        RECT  0.955 0.465 1.185 1.185 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.890 1.655 2.730 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 1.655 5.495 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.410 1.655 9.380 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.880 -0.235 10.080 0.235 ;
        RECT  9.530 -0.235 9.880 0.670 ;
        RECT  8.440 -0.235 9.530 0.235 ;
        RECT  8.090 -0.235 8.440 0.670 ;
        RECT  7.010 -0.235 8.090 0.235 ;
        RECT  6.660 -0.235 7.010 0.670 ;
        RECT  6.280 -0.235 6.660 0.235 ;
        RECT  5.930 -0.235 6.280 0.670 ;
        RECT  4.840 -0.235 5.930 0.235 ;
        RECT  4.490 -0.235 4.840 0.670 ;
        RECT  3.400 -0.235 4.490 0.235 ;
        RECT  3.050 -0.235 3.400 0.670 ;
        RECT  1.960 -0.235 3.050 0.235 ;
        RECT  1.610 -0.235 1.960 0.670 ;
        RECT  0.520 -0.235 1.610 0.235 ;
        RECT  0.170 -0.235 0.520 0.670 ;
        RECT  0.000 -0.235 0.170 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.710 3.685 10.080 4.155 ;
        RECT  2.330 2.970 2.710 4.155 ;
        RECT  1.270 3.685 2.330 4.155 ;
        RECT  0.890 2.970 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 3.055 9.160 3.285 ;
        RECT  3.345 2.475 6.280 2.705 ;
        RECT  3.115 2.475 3.345 3.330 ;
        RECT  1.905 2.475 3.115 2.705 ;
        RECT  1.675 2.475 1.905 3.330 ;
        RECT  0.465 2.475 1.675 2.710 ;
        RECT  0.235 2.475 0.465 3.330 ;
    END
END NR3D2BWP7T

MACRO NR3D3BWP7T
    CLASS CORE ;
    FOREIGN NR3D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.760 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.0610 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.195 0.480 11.425 1.180 ;
        RECT  11.195 2.380 11.425 3.295 ;
        RECT  9.985 0.900 11.195 1.180 ;
        RECT  9.130 2.380 11.195 2.680 ;
        RECT  9.755 0.480 9.985 1.180 ;
        RECT  9.130 0.900 9.755 1.180 ;
        RECT  8.545 0.900 9.130 2.680 ;
        RECT  8.315 0.480 8.545 2.680 ;
        RECT  8.230 0.900 8.315 2.680 ;
        RECT  7.105 0.900 8.230 1.180 ;
        RECT  6.875 0.480 7.105 1.180 ;
        RECT  5.665 0.900 6.875 1.180 ;
        RECT  5.435 0.480 5.665 1.180 ;
        RECT  4.225 0.900 5.435 1.180 ;
        RECT  3.995 0.480 4.225 1.180 ;
        RECT  2.785 0.900 3.995 1.180 ;
        RECT  2.555 0.480 2.785 1.180 ;
        RECT  1.345 0.900 2.555 1.180 ;
        RECT  1.115 0.480 1.345 1.180 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 2.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.425 3.630 1.655 ;
        RECT  0.700 1.425 1.540 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 2.0205 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.460 1.425 7.310 1.655 ;
        RECT  4.620 1.425 5.460 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.500 1.425 10.940 1.655 ;
        RECT  9.660 1.425 10.500 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.810 -0.235 11.760 0.235 ;
        RECT  10.410 -0.235 10.810 0.670 ;
        RECT  9.370 -0.235 10.410 0.235 ;
        RECT  8.970 -0.235 9.370 0.670 ;
        RECT  7.930 -0.235 8.970 0.235 ;
        RECT  7.530 -0.235 7.930 0.670 ;
        RECT  6.490 -0.235 7.530 0.235 ;
        RECT  6.090 -0.235 6.490 0.670 ;
        RECT  5.050 -0.235 6.090 0.235 ;
        RECT  4.650 -0.235 5.050 0.670 ;
        RECT  3.610 -0.235 4.650 0.235 ;
        RECT  3.210 -0.235 3.610 0.670 ;
        RECT  2.170 -0.235 3.210 0.235 ;
        RECT  1.770 -0.235 2.170 0.670 ;
        RECT  0.730 -0.235 1.770 0.235 ;
        RECT  0.330 -0.235 0.730 0.670 ;
        RECT  0.000 -0.235 0.330 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 3.685 11.760 4.155 ;
        RECT  3.210 2.595 3.590 4.155 ;
        RECT  2.150 3.685 3.210 4.155 ;
        RECT  1.770 3.005 2.150 4.155 ;
        RECT  0.710 3.685 1.770 4.155 ;
        RECT  0.330 2.545 0.710 4.155 ;
        RECT  0.000 3.685 0.330 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.825 3.070 10.760 3.300 ;
        RECT  7.595 2.020 7.825 3.300 ;
        RECT  4.660 3.070 7.595 3.300 ;
        RECT  4.225 2.425 7.160 2.655 ;
        RECT  3.995 2.020 4.225 3.300 ;
        RECT  2.785 2.020 3.995 2.300 ;
        RECT  2.555 2.020 2.785 3.300 ;
        RECT  1.345 2.425 2.555 2.705 ;
        RECT  1.115 2.425 1.345 3.300 ;
    END
END NR3D3BWP7T

MACRO NR3D4BWP7T
    CLASS CORE ;
    FOREIGN NR3D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 6.5964 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.535 2.505 15.775 3.370 ;
        RECT  15.540 0.515 15.770 1.250 ;
        RECT  14.330 0.900 15.540 1.250 ;
        RECT  12.945 2.505 15.535 2.855 ;
        RECT  14.100 0.515 14.330 1.250 ;
        RECT  12.890 0.900 14.100 1.250 ;
        RECT  12.600 2.100 12.945 2.855 ;
        RECT  12.660 0.515 12.890 1.250 ;
        RECT  11.930 0.900 12.660 1.250 ;
        RECT  11.930 2.100 12.600 2.415 ;
        RECT  11.505 0.900 11.930 2.415 ;
        RECT  11.450 0.900 11.505 2.855 ;
        RECT  11.220 0.515 11.450 2.855 ;
        RECT  11.030 0.900 11.220 2.855 ;
        RECT  10.010 0.900 11.030 1.250 ;
        RECT  9.780 0.515 10.010 1.250 ;
        RECT  8.570 0.900 9.780 1.250 ;
        RECT  8.340 0.515 8.570 1.250 ;
        RECT  7.130 0.900 8.340 1.250 ;
        RECT  6.900 0.515 7.130 1.250 ;
        RECT  5.690 0.900 6.900 1.250 ;
        RECT  5.460 0.515 5.690 1.250 ;
        RECT  4.250 0.900 5.460 1.250 ;
        RECT  4.020 0.515 4.250 1.250 ;
        RECT  2.810 0.900 4.020 1.250 ;
        RECT  2.580 0.515 2.810 1.250 ;
        RECT  1.370 0.900 2.580 1.250 ;
        RECT  1.140 0.515 1.370 1.250 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 2.6910 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.480 5.100 1.710 ;
        RECT  0.700 1.480 1.540 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 2.7342 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.700 1.480 10.175 1.710 ;
        RECT  7.420 1.480 7.700 2.150 ;
        RECT  6.580 1.480 7.420 1.710 ;
        RECT  6.300 1.480 6.580 2.150 ;
        RECT  6.075 1.480 6.300 1.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.6910 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.700 1.480 15.540 2.150 ;
        RECT  12.185 1.480 14.700 1.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.135 -0.235 16.240 0.235 ;
        RECT  14.750 -0.235 15.135 0.670 ;
        RECT  13.695 -0.235 14.750 0.235 ;
        RECT  13.310 -0.235 13.695 0.670 ;
        RECT  12.255 -0.235 13.310 0.235 ;
        RECT  11.870 -0.235 12.255 0.670 ;
        RECT  10.835 -0.235 11.870 0.235 ;
        RECT  10.395 -0.235 10.835 0.670 ;
        RECT  9.375 -0.235 10.395 0.235 ;
        RECT  8.990 -0.235 9.375 0.670 ;
        RECT  7.935 -0.235 8.990 0.235 ;
        RECT  7.550 -0.235 7.935 0.670 ;
        RECT  6.495 -0.235 7.550 0.235 ;
        RECT  6.110 -0.235 6.495 0.670 ;
        RECT  5.055 -0.235 6.110 0.235 ;
        RECT  4.670 -0.235 5.055 0.670 ;
        RECT  3.615 -0.235 4.670 0.235 ;
        RECT  3.230 -0.235 3.615 0.670 ;
        RECT  2.175 -0.235 3.230 0.235 ;
        RECT  1.790 -0.235 2.175 0.670 ;
        RECT  0.735 -0.235 1.790 0.235 ;
        RECT  0.350 -0.235 0.735 0.670 ;
        RECT  0.000 -0.235 0.350 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.050 3.685 16.240 4.155 ;
        RECT  4.670 2.620 5.050 4.155 ;
        RECT  3.610 3.685 4.670 4.155 ;
        RECT  3.230 2.620 3.610 4.155 ;
        RECT  2.170 3.685 3.230 4.155 ;
        RECT  1.790 3.125 2.170 4.155 ;
        RECT  0.730 3.685 1.790 4.155 ;
        RECT  0.350 2.560 0.730 4.155 ;
        RECT  0.000 3.685 0.350 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.535 2.505 15.775 3.370 ;
        RECT  15.540 0.515 15.770 1.250 ;
        RECT  14.330 0.900 15.540 1.250 ;
        RECT  12.945 2.505 15.535 2.855 ;
        RECT  14.100 0.515 14.330 1.250 ;
        RECT  12.890 0.900 14.100 1.250 ;
        RECT  12.600 2.100 12.945 2.855 ;
        RECT  12.660 0.515 12.890 1.250 ;
        RECT  12.130 0.900 12.660 1.250 ;
        RECT  12.130 2.100 12.600 2.415 ;
        RECT  10.010 0.900 10.830 1.250 ;
        RECT  9.780 0.515 10.010 1.250 ;
        RECT  8.570 0.900 9.780 1.250 ;
        RECT  8.340 0.515 8.570 1.250 ;
        RECT  7.130 0.900 8.340 1.250 ;
        RECT  6.900 0.515 7.130 1.250 ;
        RECT  5.690 0.900 6.900 1.250 ;
        RECT  5.460 0.515 5.690 1.250 ;
        RECT  4.250 0.900 5.460 1.250 ;
        RECT  4.020 0.515 4.250 1.250 ;
        RECT  2.810 0.900 4.020 1.250 ;
        RECT  2.580 0.515 2.810 1.250 ;
        RECT  1.370 0.900 2.580 1.250 ;
        RECT  1.140 0.515 1.370 1.250 ;
        RECT  12.225 3.135 15.105 3.365 ;
        RECT  11.885 2.660 12.225 3.365 ;
        RECT  10.730 3.135 11.885 3.365 ;
        RECT  10.500 2.140 10.730 3.365 ;
        RECT  9.300 3.135 10.500 3.365 ;
        RECT  9.780 2.045 10.010 2.860 ;
        RECT  8.570 2.045 9.780 2.335 ;
        RECT  9.050 2.585 9.300 3.365 ;
        RECT  6.125 3.135 9.050 3.365 ;
        RECT  8.340 2.045 8.570 2.860 ;
        RECT  7.130 2.570 8.340 2.860 ;
        RECT  6.900 2.100 7.130 2.860 ;
        RECT  5.690 2.555 6.900 2.860 ;
        RECT  5.460 2.030 5.690 3.310 ;
        RECT  4.250 2.030 5.460 2.330 ;
        RECT  4.020 2.030 4.250 3.310 ;
        RECT  2.810 2.045 4.020 2.330 ;
        RECT  2.580 2.045 2.810 3.360 ;
        RECT  1.370 2.570 2.580 2.855 ;
        RECT  1.140 2.570 1.370 3.380 ;
    END
END NR3D4BWP7T

MACRO NR4D0BWP7T
    CLASS CORE ;
    FOREIGN NR4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2051 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.880 2.245 3.110 3.455 ;
        RECT  1.030 3.225 2.880 3.455 ;
        RECT  0.980 0.855 2.580 1.085 ;
        RECT  0.980 2.755 1.030 3.455 ;
        RECT  0.800 0.855 0.980 3.455 ;
        RECT  0.700 0.855 0.800 2.985 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.580 0.450 2.710 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.580 1.540 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.580 2.200 1.920 ;
        RECT  1.820 1.580 2.100 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.650 3.220 1.670 ;
        RECT  2.585 1.440 2.940 1.670 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.525 -0.235 3.360 0.235 ;
        RECT  0.470 -0.235 0.525 0.420 ;
        RECT  0.145 -0.235 0.470 1.140 ;
        RECT  0.000 -0.235 0.145 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 3.685 3.360 4.155 ;
        RECT  0.155 3.160 0.535 4.155 ;
        RECT  0.000 3.685 0.155 4.155 ;
        END
    END VDD
END NR4D0BWP7T

MACRO NR4D1BWP7T
    CLASS CORE ;
    FOREIGN NR4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8198 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.355 0.800 3.980 1.030 ;
        RECT  0.355 2.380 1.780 2.660 ;
        RECT  0.125 0.800 0.355 2.660 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.770 4.900 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.260 5.460 1.940 ;
        RECT  3.305 1.260 5.150 1.540 ;
        RECT  3.075 1.260 3.305 1.825 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.260 2.660 2.150 ;
        RECT  0.815 1.260 2.380 1.540 ;
        RECT  0.585 1.260 0.815 2.065 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 1.770 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.700 -0.235 5.600 0.235 ;
        RECT  4.340 -0.235 4.700 0.845 ;
        RECT  3.230 -0.235 4.340 0.235 ;
        RECT  2.855 -0.235 3.230 0.570 ;
        RECT  1.710 -0.235 2.855 0.235 ;
        RECT  1.345 -0.235 1.710 0.570 ;
        RECT  0.000 -0.235 1.345 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.290 3.685 5.600 4.155 ;
        RECT  3.890 2.940 4.290 4.155 ;
        RECT  0.000 3.685 3.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.135 2.410 5.365 3.400 ;
        RECT  3.495 2.410 5.135 2.640 ;
        RECT  3.265 2.410 3.495 3.120 ;
        RECT  0.180 2.890 3.265 3.120 ;
    END
END NR4D1BWP7T

MACRO NR4D2BWP7T
    CLASS CORE ;
    FOREIGN NR4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 4.1796 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.415 0.465 12.645 1.180 ;
        RECT  11.205 0.900 12.415 1.180 ;
        RECT  10.250 2.500 11.980 2.780 ;
        RECT  10.975 0.465 11.205 1.180 ;
        RECT  10.250 0.900 10.975 1.180 ;
        RECT  10.000 0.900 10.250 2.780 ;
        RECT  9.765 0.900 10.000 2.430 ;
        RECT  9.535 0.465 9.765 2.430 ;
        RECT  9.350 0.900 9.535 2.430 ;
        RECT  8.325 0.900 9.350 1.180 ;
        RECT  8.095 0.465 8.325 1.180 ;
        RECT  6.940 0.900 8.095 1.180 ;
        RECT  5.940 0.480 6.940 1.180 ;
        RECT  4.785 0.900 5.940 1.180 ;
        RECT  4.555 0.465 4.785 1.180 ;
        RECT  3.345 0.900 4.555 1.180 ;
        RECT  3.115 0.465 3.345 1.180 ;
        RECT  1.905 0.900 3.115 1.180 ;
        RECT  1.675 0.465 1.905 1.180 ;
        RECT  0.465 0.900 1.675 1.180 ;
        RECT  0.235 0.465 0.465 1.180 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.410 2.580 1.640 ;
        RECT  1.260 1.410 2.110 2.150 ;
        RECT  0.730 1.410 1.260 1.640 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.460 1.410 5.630 1.640 ;
        RECT  4.620 1.410 5.460 2.150 ;
        RECT  3.780 1.410 4.620 1.640 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 1.410 9.095 1.640 ;
        RECT  7.865 1.410 8.820 2.150 ;
        RECT  7.245 1.410 7.865 1.640 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.3464 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.655 1.410 11.620 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.030 -0.235 12.880 0.235 ;
        RECT  11.630 -0.235 12.030 0.670 ;
        RECT  10.590 -0.235 11.630 0.235 ;
        RECT  10.190 -0.235 10.590 0.670 ;
        RECT  9.150 -0.235 10.190 0.235 ;
        RECT  8.750 -0.235 9.150 0.670 ;
        RECT  7.710 -0.235 8.750 0.235 ;
        RECT  7.310 -0.235 7.710 0.670 ;
        RECT  5.610 -0.235 7.310 0.235 ;
        RECT  5.210 -0.235 5.610 0.670 ;
        RECT  4.170 -0.235 5.210 0.235 ;
        RECT  3.770 -0.235 4.170 0.670 ;
        RECT  2.730 -0.235 3.770 0.235 ;
        RECT  2.330 -0.235 2.730 0.670 ;
        RECT  1.290 -0.235 2.330 0.235 ;
        RECT  0.890 -0.235 1.290 0.670 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.710 3.685 12.880 4.155 ;
        RECT  2.330 3.005 2.710 4.155 ;
        RECT  1.270 3.685 2.330 4.155 ;
        RECT  0.890 3.005 1.270 4.155 ;
        RECT  0.000 3.685 0.890 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.415 2.535 12.645 3.455 ;
        RECT  6.600 3.225 12.415 3.455 ;
        RECT  6.370 2.765 9.100 2.995 ;
        RECT  6.140 2.765 6.370 3.330 ;
        RECT  5.930 2.305 6.320 2.535 ;
        RECT  3.780 3.100 6.140 3.330 ;
        RECT  5.700 2.305 5.930 2.620 ;
        RECT  3.345 2.380 5.700 2.620 ;
        RECT  3.115 2.380 3.345 3.255 ;
        RECT  1.905 2.380 3.115 2.620 ;
        RECT  1.675 2.380 1.905 3.360 ;
        RECT  0.465 2.380 1.675 2.620 ;
        RECT  0.235 2.380 0.465 3.360 ;
    END
END NR4D2BWP7T

MACRO NR4D3BWP7T
    CLASS CORE ;
    FOREIGN NR4D3BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 6.1122 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.845 0.515 15.075 1.200 ;
        RECT  14.845 2.460 15.075 3.360 ;
        RECT  13.635 0.900 14.845 1.200 ;
        RECT  12.490 2.460 14.845 2.780 ;
        RECT  13.405 0.515 13.635 1.200 ;
        RECT  12.490 0.900 13.405 1.200 ;
        RECT  12.195 0.900 12.490 2.780 ;
        RECT  11.965 0.515 12.195 2.780 ;
        RECT  11.590 0.900 11.965 2.780 ;
        RECT  10.755 0.900 11.590 1.200 ;
        RECT  10.525 0.515 10.755 1.200 ;
        RECT  9.315 0.900 10.525 1.200 ;
        RECT  9.085 0.515 9.315 1.200 ;
        RECT  7.875 0.900 9.085 1.200 ;
        RECT  7.645 0.515 7.875 1.200 ;
        RECT  6.435 0.900 7.645 1.200 ;
        RECT  6.205 0.515 6.435 1.200 ;
        RECT  4.995 0.900 6.205 1.200 ;
        RECT  4.765 0.515 4.995 1.200 ;
        RECT  3.555 0.900 4.765 1.200 ;
        RECT  3.325 0.515 3.555 1.200 ;
        RECT  2.115 0.900 3.325 1.200 ;
        RECT  1.885 0.515 2.115 1.200 ;
        RECT  0.675 0.900 1.885 1.200 ;
        RECT  0.445 0.515 0.675 1.200 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 2.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.430 3.685 1.660 ;
        RECT  1.820 1.430 2.660 2.150 ;
        RECT  0.995 1.430 1.820 1.660 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 2.0205 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.580 1.430 7.280 1.660 ;
        RECT  5.740 1.430 6.580 2.150 ;
        RECT  4.590 1.430 5.740 1.660 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 2.0205 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.940 1.430 10.570 1.660 ;
        RECT  9.100 1.430 9.940 2.150 ;
        RECT  8.350 1.430 9.100 1.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.0196 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.430 14.140 2.150 ;
        RECT  12.860 1.430 13.020 1.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.440 -0.235 15.680 0.235 ;
        RECT  14.060 -0.235 14.440 0.670 ;
        RECT  13.000 -0.235 14.060 0.235 ;
        RECT  12.620 -0.235 13.000 0.670 ;
        RECT  11.560 -0.235 12.620 0.235 ;
        RECT  11.180 -0.235 11.560 0.670 ;
        RECT  10.120 -0.235 11.180 0.235 ;
        RECT  9.740 -0.235 10.120 0.670 ;
        RECT  8.680 -0.235 9.740 0.235 ;
        RECT  8.300 -0.235 8.680 0.670 ;
        RECT  7.240 -0.235 8.300 0.235 ;
        RECT  6.860 -0.235 7.240 0.670 ;
        RECT  5.800 -0.235 6.860 0.235 ;
        RECT  5.420 -0.235 5.800 0.670 ;
        RECT  4.360 -0.235 5.420 0.235 ;
        RECT  3.980 -0.235 4.360 0.670 ;
        RECT  2.920 -0.235 3.980 0.235 ;
        RECT  2.540 -0.235 2.920 0.670 ;
        RECT  1.480 -0.235 2.540 0.235 ;
        RECT  1.100 -0.235 1.480 0.670 ;
        RECT  0.000 -0.235 1.100 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.640 3.685 15.680 4.155 ;
        RECT  3.260 3.005 3.640 4.155 ;
        RECT  2.200 3.685 3.260 4.155 ;
        RECT  1.820 3.005 2.200 4.155 ;
        RECT  0.760 3.685 1.820 4.155 ;
        RECT  0.380 2.635 0.760 4.155 ;
        RECT  0.000 3.685 0.380 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.845 0.515 15.075 1.200 ;
        RECT  14.845 2.460 15.075 3.360 ;
        RECT  13.635 0.900 14.845 1.200 ;
        RECT  12.690 2.460 14.845 2.780 ;
        RECT  13.405 0.515 13.635 1.200 ;
        RECT  12.690 0.900 13.405 1.200 ;
        RECT  10.755 0.900 11.390 1.200 ;
        RECT  10.525 0.515 10.755 1.200 ;
        RECT  9.315 0.900 10.525 1.200 ;
        RECT  9.085 0.515 9.315 1.200 ;
        RECT  7.875 0.900 9.085 1.200 ;
        RECT  7.645 0.515 7.875 1.200 ;
        RECT  6.435 0.900 7.645 1.200 ;
        RECT  6.205 0.515 6.435 1.200 ;
        RECT  4.995 0.900 6.205 1.200 ;
        RECT  4.765 0.515 4.995 1.200 ;
        RECT  3.555 0.900 4.765 1.200 ;
        RECT  3.325 0.515 3.555 1.200 ;
        RECT  2.115 0.900 3.325 1.200 ;
        RECT  1.885 0.515 2.115 1.200 ;
        RECT  0.675 0.900 1.885 1.200 ;
        RECT  0.445 0.515 0.675 1.200 ;
        RECT  8.310 3.055 14.410 3.285 ;
        RECT  10.525 1.975 10.755 2.785 ;
        RECT  7.875 2.555 10.525 2.785 ;
        RECT  7.645 2.010 7.875 3.290 ;
        RECT  4.710 2.555 7.645 2.785 ;
        RECT  4.275 3.070 7.210 3.300 ;
        RECT  4.045 2.020 4.275 3.300 ;
        RECT  2.835 2.490 4.045 2.730 ;
        RECT  2.605 2.490 2.835 3.360 ;
        RECT  1.395 2.490 2.605 2.730 ;
        RECT  1.165 2.490 1.395 3.360 ;
    END
END NR4D3BWP7T

MACRO NR4D4BWP7T
    CLASS CORE ;
    FOREIGN NR4D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 7.6384 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.600 2.380 20.830 3.200 ;
        RECT  16.970 2.380 20.600 2.730 ;
        RECT  19.880 0.525 20.110 1.250 ;
        RECT  18.670 0.900 19.880 1.250 ;
        RECT  18.440 0.525 18.670 1.250 ;
        RECT  17.230 0.900 18.440 1.250 ;
        RECT  17.000 0.525 17.230 1.250 ;
        RECT  16.970 0.900 17.000 1.250 ;
        RECT  16.070 0.900 16.970 2.730 ;
        RECT  15.790 0.900 16.070 1.250 ;
        RECT  15.560 0.525 15.790 1.250 ;
        RECT  14.350 0.900 15.560 1.250 ;
        RECT  14.120 0.525 14.350 1.250 ;
        RECT  12.910 0.900 14.120 1.250 ;
        RECT  12.680 0.525 12.910 1.250 ;
        RECT  11.470 0.900 12.680 1.250 ;
        RECT  11.240 0.525 11.470 1.250 ;
        RECT  10.030 0.900 11.240 1.250 ;
        RECT  9.800 0.525 10.030 1.250 ;
        RECT  8.590 0.900 9.800 1.250 ;
        RECT  8.360 0.525 8.590 1.250 ;
        RECT  7.150 0.900 8.360 1.250 ;
        RECT  6.920 0.525 7.150 1.250 ;
        RECT  5.710 0.900 6.920 1.250 ;
        RECT  5.480 0.525 5.710 1.250 ;
        RECT  4.270 0.900 5.480 1.250 ;
        RECT  4.040 0.525 4.270 1.250 ;
        RECT  2.830 0.900 4.040 1.250 ;
        RECT  2.600 0.525 2.830 1.250 ;
        RECT  1.390 0.900 2.600 1.250 ;
        RECT  1.160 0.525 1.390 1.250 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 2.6910 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.480 5.060 1.710 ;
        RECT  0.700 1.480 1.540 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 2.7342 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.580 1.480 10.285 1.710 ;
        RECT  5.740 1.480 6.580 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 2.7342 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.140 1.480 15.095 2.150 ;
        RECT  10.995 1.480 14.140 1.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 2.6910 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.340 1.480 20.395 1.710 ;
        RECT  17.500 1.480 18.340 2.150 ;
        RECT  17.235 1.480 17.500 1.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  20.920 -0.235 21.280 0.235 ;
        RECT  20.530 -0.235 20.920 0.745 ;
        RECT  19.480 -0.235 20.530 0.235 ;
        RECT  19.090 -0.235 19.480 0.670 ;
        RECT  18.040 -0.235 19.090 0.235 ;
        RECT  17.650 -0.235 18.040 0.670 ;
        RECT  16.600 -0.235 17.650 0.235 ;
        RECT  16.210 -0.235 16.600 0.670 ;
        RECT  15.160 -0.235 16.210 0.235 ;
        RECT  14.770 -0.235 15.160 0.670 ;
        RECT  13.720 -0.235 14.770 0.235 ;
        RECT  13.330 -0.235 13.720 0.670 ;
        RECT  12.280 -0.235 13.330 0.235 ;
        RECT  11.890 -0.235 12.280 0.670 ;
        RECT  10.830 -0.235 11.890 0.235 ;
        RECT  10.415 -0.235 10.830 0.670 ;
        RECT  9.400 -0.235 10.415 0.235 ;
        RECT  9.010 -0.235 9.400 0.670 ;
        RECT  7.960 -0.235 9.010 0.235 ;
        RECT  7.570 -0.235 7.960 0.670 ;
        RECT  6.520 -0.235 7.570 0.235 ;
        RECT  6.130 -0.235 6.520 0.670 ;
        RECT  5.080 -0.235 6.130 0.235 ;
        RECT  4.690 -0.235 5.080 0.670 ;
        RECT  3.640 -0.235 4.690 0.235 ;
        RECT  3.250 -0.235 3.640 0.670 ;
        RECT  2.200 -0.235 3.250 0.235 ;
        RECT  1.810 -0.235 2.200 0.670 ;
        RECT  0.755 -0.235 1.810 0.235 ;
        RECT  0.365 -0.235 0.755 0.770 ;
        RECT  0.000 -0.235 0.365 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.070 3.685 21.280 4.155 ;
        RECT  4.690 3.080 5.070 4.155 ;
        RECT  3.630 3.685 4.690 4.155 ;
        RECT  3.250 2.630 3.630 4.155 ;
        RECT  2.190 3.685 3.250 4.155 ;
        RECT  1.810 3.080 2.190 4.155 ;
        RECT  0.745 3.685 1.810 4.155 ;
        RECT  0.360 2.610 0.745 4.155 ;
        RECT  0.000 3.685 0.360 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.600 2.380 20.830 3.200 ;
        RECT  17.170 2.380 20.600 2.730 ;
        RECT  19.880 0.525 20.110 1.250 ;
        RECT  18.670 0.900 19.880 1.250 ;
        RECT  18.440 0.525 18.670 1.250 ;
        RECT  17.230 0.900 18.440 1.250 ;
        RECT  17.170 0.525 17.230 1.250 ;
        RECT  15.790 0.900 15.870 1.250 ;
        RECT  15.560 0.525 15.790 1.250 ;
        RECT  14.350 0.900 15.560 1.250 ;
        RECT  14.120 0.525 14.350 1.250 ;
        RECT  12.910 0.900 14.120 1.250 ;
        RECT  12.680 0.525 12.910 1.250 ;
        RECT  11.470 0.900 12.680 1.250 ;
        RECT  11.240 0.525 11.470 1.250 ;
        RECT  10.030 0.900 11.240 1.250 ;
        RECT  9.800 0.525 10.030 1.250 ;
        RECT  8.590 0.900 9.800 1.250 ;
        RECT  8.360 0.525 8.590 1.250 ;
        RECT  7.150 0.900 8.360 1.250 ;
        RECT  6.920 0.525 7.150 1.250 ;
        RECT  5.710 0.900 6.920 1.250 ;
        RECT  5.480 0.525 5.710 1.250 ;
        RECT  4.270 0.900 5.480 1.250 ;
        RECT  4.040 0.525 4.270 1.250 ;
        RECT  2.830 0.900 4.040 1.250 ;
        RECT  2.600 0.525 2.830 1.250 ;
        RECT  1.390 0.900 2.600 1.250 ;
        RECT  1.160 0.525 1.390 1.250 ;
        RECT  15.790 3.100 20.165 3.380 ;
        RECT  15.560 2.080 15.790 3.380 ;
        RECT  11.185 3.100 15.560 3.380 ;
        RECT  10.750 2.435 15.125 2.695 ;
        RECT  10.520 2.435 10.750 3.205 ;
        RECT  6.065 2.435 10.520 2.695 ;
        RECT  5.710 3.090 10.085 3.370 ;
        RECT  5.480 2.560 5.710 3.370 ;
        RECT  4.270 2.560 5.480 2.850 ;
        RECT  4.040 2.080 4.270 3.370 ;
        RECT  2.830 2.080 4.040 2.370 ;
        RECT  2.600 2.080 2.830 3.360 ;
        RECT  1.385 2.560 2.600 2.850 ;
        RECT  1.155 2.560 1.385 3.370 ;
    END
END NR4D4BWP7T

MACRO OA211D0BWP7T
    CLASS CORE ;
    FOREIGN OA211D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5962 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.520 4.340 3.345 ;
        RECT  3.960 0.520 4.060 0.750 ;
        RECT  3.785 3.115 4.060 3.345 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.010 2.330 1.485 2.560 ;
        RECT  0.700 1.210 1.010 2.560 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.570 1.630 2.070 1.860 ;
        RECT  1.260 0.650 1.570 1.860 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.210 3.225 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 -0.235 4.480 0.235 ;
        RECT  3.235 -0.235 3.615 0.750 ;
        RECT  0.620 -0.235 3.235 0.235 ;
        RECT  0.180 -0.235 0.620 0.670 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 3.685 4.480 4.155 ;
        RECT  2.920 3.115 3.300 4.155 ;
        RECT  1.290 3.685 2.920 4.155 ;
        RECT  0.905 3.250 1.290 4.155 ;
        RECT  0.000 3.685 0.905 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.560 1.625 3.790 2.885 ;
        RECT  2.600 2.645 3.560 2.885 ;
        RECT  2.370 0.815 2.600 3.020 ;
        RECT  1.970 0.815 2.370 1.045 ;
        RECT  1.945 2.790 2.370 3.020 ;
        RECT  1.680 2.790 1.945 3.390 ;
        RECT  0.485 2.790 1.680 3.020 ;
        RECT  0.255 2.790 0.485 3.370 ;
    END
END OA211D0BWP7T

MACRO OA211D1BWP7T
    CLASS CORE ;
    FOREIGN OA211D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.560 0.470 4.900 3.300 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.715 0.980 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.210 1.540 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.715 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.905 1.715 3.785 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 -0.235 5.040 0.235 ;
        RECT  3.760 -0.235 4.140 0.790 ;
        RECT  0.600 -0.235 3.760 0.235 ;
        RECT  0.220 -0.235 0.600 1.215 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.150 3.685 5.040 4.155 ;
        RECT  3.770 2.995 4.150 4.155 ;
        RECT  3.350 3.685 3.770 4.155 ;
        RECT  2.970 2.995 3.350 4.155 ;
        RECT  1.310 3.685 2.970 4.155 ;
        RECT  0.930 2.995 1.310 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.040 1.020 4.270 2.730 ;
        RECT  2.265 1.020 4.040 1.250 ;
        RECT  1.945 2.450 4.040 2.730 ;
        RECT  1.540 0.535 3.325 0.765 ;
        RECT  1.715 2.450 1.945 3.320 ;
        RECT  0.505 2.450 1.715 2.730 ;
        RECT  0.275 2.450 0.505 3.320 ;
    END
END OA211D1BWP7T

MACRO OA211D2BWP7T
    CLASS CORE ;
    FOREIGN OA211D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.645 1.210 4.900 2.235 ;
        RECT  4.620 0.465 4.645 3.370 ;
        RECT  4.415 0.465 4.620 1.440 ;
        RECT  4.415 2.005 4.620 3.370 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 1.210 1.560 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.695 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.625 3.220 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.365 -0.235 5.600 0.235 ;
        RECT  5.135 -0.235 5.365 1.245 ;
        RECT  3.980 -0.235 5.135 0.235 ;
        RECT  3.640 -0.235 3.980 0.670 ;
        RECT  0.465 -0.235 3.640 0.235 ;
        RECT  0.235 -0.235 0.465 1.230 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.365 3.685 5.600 4.155 ;
        RECT  5.135 2.475 5.365 4.155 ;
        RECT  3.940 3.685 5.135 4.155 ;
        RECT  3.600 3.455 3.940 4.155 ;
        RECT  3.200 3.685 3.600 4.155 ;
        RECT  2.860 3.455 3.200 4.155 ;
        RECT  1.265 3.685 2.860 4.155 ;
        RECT  0.885 2.900 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.955 0.925 4.185 3.225 ;
        RECT  2.100 0.925 3.955 1.155 ;
        RECT  1.905 2.985 3.955 3.225 ;
        RECT  1.375 0.465 3.160 0.695 ;
        RECT  1.675 2.380 1.905 3.225 ;
        RECT  0.465 2.380 1.675 2.610 ;
        RECT  0.235 2.380 0.465 3.320 ;
    END
END OA211D2BWP7T

MACRO OA21D0BWP7T
    CLASS CORE ;
    FOREIGN OA21D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 0.570 3.220 3.175 ;
        RECT  2.840 0.570 2.940 0.800 ;
        RECT  2.840 2.945 2.940 3.175 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.660 1.590 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.600 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.480 -0.235 3.360 0.235 ;
        RECT  2.100 -0.235 2.480 0.820 ;
        RECT  0.000 -0.235 2.100 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.430 3.685 3.360 4.155 ;
        RECT  2.070 3.455 2.430 4.155 ;
        RECT  0.520 3.685 2.070 4.155 ;
        RECT  0.180 3.455 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.480 1.855 2.710 2.740 ;
        RECT  1.025 2.510 2.480 2.740 ;
        RECT  0.795 0.830 1.025 2.740 ;
    END
END OA21D0BWP7T

MACRO OA21D1BWP7T
    CLASS CORE ;
    FOREIGN OA21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 1.210 3.780 2.710 ;
        RECT  3.685 1.210 3.695 3.345 ;
        RECT  3.500 0.465 3.685 3.345 ;
        RECT  3.455 0.465 3.500 1.470 ;
        RECT  3.455 2.375 3.500 3.345 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.210 2.660 2.150 ;
        RECT  2.330 1.680 2.380 2.020 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.620 0.465 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 2.150 ;
        RECT  1.530 1.735 1.820 1.965 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 -0.235 3.920 0.235 ;
        RECT  2.680 -0.235 3.020 0.730 ;
        RECT  0.000 -0.235 2.680 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.050 3.685 3.920 4.155 ;
        RECT  2.670 3.025 3.050 4.155 ;
        RECT  0.600 3.685 2.670 4.155 ;
        RECT  0.220 3.025 0.600 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.185 1.650 3.250 2.045 ;
        RECT  3.020 1.650 3.185 2.670 ;
        RECT  2.955 1.815 3.020 2.670 ;
        RECT  2.180 2.430 2.955 2.670 ;
        RECT  1.950 0.465 2.180 0.960 ;
        RECT  1.950 2.430 2.180 3.345 ;
        RECT  0.505 0.465 1.950 0.705 ;
        RECT  1.230 2.430 1.950 2.670 ;
        RECT  0.990 0.965 1.230 2.670 ;
        RECT  0.275 0.465 0.505 0.960 ;
    END
END OA21D1BWP7T

MACRO OA21D2BWP7T
    CLASS CORE ;
    FOREIGN OA21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.475 3.780 3.175 ;
        RECT  3.230 0.475 3.500 0.705 ;
        RECT  3.240 2.945 3.500 3.175 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.735 2.660 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.725 0.465 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.560 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 -0.235 4.480 0.235 ;
        RECT  4.010 -0.235 4.245 1.325 ;
        RECT  2.860 -0.235 4.010 0.235 ;
        RECT  2.520 -0.235 2.860 0.670 ;
        RECT  0.000 -0.235 2.520 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 3.685 4.480 4.155 ;
        RECT  4.015 2.245 4.245 4.155 ;
        RECT  2.880 3.685 4.015 4.155 ;
        RECT  2.500 2.935 2.880 4.155 ;
        RECT  0.600 3.685 2.500 4.155 ;
        RECT  0.220 3.025 0.600 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.040 0.935 3.270 2.670 ;
        RECT  0.915 0.935 3.040 1.165 ;
        RECT  2.005 2.430 3.040 2.670 ;
        RECT  0.505 0.465 2.070 0.695 ;
        RECT  1.775 2.430 2.005 3.330 ;
        RECT  0.275 0.465 0.505 1.275 ;
    END
END OA21D2BWP7T

MACRO OA221D0BWP7T
    CLASS CORE ;
    FOREIGN OA221D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 0.465 4.900 3.410 ;
        RECT  4.440 0.465 4.620 0.695 ;
        RECT  4.575 3.070 4.620 3.410 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 2.380 3.830 2.660 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.820 3.270 2.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.450 2.380 2.400 2.660 ;
        RECT  0.220 1.015 0.450 2.660 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.675 2.100 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.070 -0.235 5.040 0.235 ;
        RECT  3.690 -0.235 4.070 0.685 ;
        RECT  0.000 -0.235 3.690 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.115 3.685 5.040 4.155 ;
        RECT  3.745 3.455 4.115 4.155 ;
        RECT  1.965 3.685 3.745 4.155 ;
        RECT  1.625 3.455 1.965 4.155 ;
        RECT  0.000 3.685 1.625 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.095 0.925 4.325 3.225 ;
        RECT  1.540 0.925 4.095 1.155 ;
        RECT  0.200 2.995 4.095 3.225 ;
        RECT  0.190 0.465 3.340 0.695 ;
    END
END OA221D0BWP7T

MACRO OA221D1BWP7T
    CLASS CORE ;
    FOREIGN OA221D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 0.465 5.460 3.230 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4005 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.720 4.350 2.150 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.680 2.115 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4005 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.735 3.220 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.680 1.540 2.710 ;
        RECT  1.185 1.680 1.260 2.040 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.715 -0.235 5.600 0.235 ;
        RECT  4.335 -0.235 4.715 1.205 ;
        RECT  0.000 -0.235 4.335 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.700 3.685 5.600 4.155 ;
        RECT  4.360 2.885 4.700 4.155 ;
        RECT  3.240 3.685 4.360 4.155 ;
        RECT  2.900 2.940 3.240 4.155 ;
        RECT  0.485 3.685 2.900 4.155 ;
        RECT  0.255 2.940 0.485 4.155 ;
        RECT  0.000 3.685 0.255 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.655 1.680 4.885 2.610 ;
        RECT  3.925 2.380 4.655 2.610 ;
        RECT  2.340 0.465 3.980 0.695 ;
        RECT  3.695 2.380 3.925 3.390 ;
        RECT  2.575 2.380 3.695 2.610 ;
        RECT  1.905 1.140 3.445 1.370 ;
        RECT  2.345 2.380 2.575 3.170 ;
        RECT  0.955 2.940 2.345 3.170 ;
        RECT  1.675 0.465 1.905 1.370 ;
        RECT  0.180 0.465 1.675 0.695 ;
        RECT  0.955 1.020 1.240 1.250 ;
        RECT  0.715 1.020 0.955 3.170 ;
    END
END OA221D1BWP7T

MACRO OA221D2BWP7T
    CLASS CORE ;
    FOREIGN OA221D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.7301 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.170 6.020 2.420 ;
        RECT  5.630 1.170 5.740 1.430 ;
        RECT  5.630 2.180 5.740 2.420 ;
        RECT  5.400 0.465 5.630 1.430 ;
        RECT  5.400 2.180 5.630 3.340 ;
        END
    END Z
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.400 2.150 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.590 3.780 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.695 3.220 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.140 1.735 2.100 2.190 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 -0.235 6.720 0.235 ;
        RECT  6.255 -0.235 6.485 1.280 ;
        RECT  4.895 -0.235 6.255 0.235 ;
        RECT  4.515 -0.235 4.895 0.945 ;
        RECT  0.000 -0.235 4.515 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 3.685 6.720 4.155 ;
        RECT  6.255 2.195 6.485 4.155 ;
        RECT  4.765 3.685 6.255 4.155 ;
        RECT  4.535 2.850 4.765 4.155 ;
        RECT  2.735 3.685 4.535 4.155 ;
        RECT  2.355 2.950 2.735 4.155 ;
        RECT  0.560 3.685 2.355 4.155 ;
        RECT  0.180 2.950 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.945 1.695 5.480 1.925 ;
        RECT  4.690 1.695 4.945 2.610 ;
        RECT  4.245 2.380 4.690 2.610 ;
        RECT  4.010 2.380 4.245 3.245 ;
        RECT  3.855 0.465 4.085 0.975 ;
        RECT  3.240 3.015 4.010 3.245 ;
        RECT  2.360 0.465 3.855 0.695 ;
        RECT  1.905 0.925 3.420 1.155 ;
        RECT  3.010 2.440 3.240 3.245 ;
        RECT  1.905 2.440 3.010 2.670 ;
        RECT  1.675 0.465 1.905 1.310 ;
        RECT  1.675 2.440 1.905 3.300 ;
        RECT  0.465 0.465 1.675 0.695 ;
        RECT  0.910 2.440 1.675 2.670 ;
        RECT  0.910 0.925 1.240 1.155 ;
        RECT  0.680 0.925 0.910 2.670 ;
        RECT  0.235 0.465 0.465 0.820 ;
    END
END OA221D2BWP7T

MACRO OA222D0BWP7T
    CLASS CORE ;
    FOREIGN OA222D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 0.980 6.020 3.355 ;
        RECT  5.640 0.980 5.740 1.210 ;
        RECT  5.640 3.125 5.740 3.355 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 1.730 1.540 2.710 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.730 2.145 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.705 4.900 2.710 ;
        RECT  2.530 2.445 4.620 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.765 3.240 2.190 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 4.340 2.195 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 -0.235 6.160 0.235 ;
        RECT  5.695 -0.235 5.925 0.540 ;
        RECT  1.270 -0.235 5.695 0.235 ;
        RECT  0.890 -0.235 1.270 0.930 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.235 3.685 6.160 4.155 ;
        RECT  4.865 3.455 5.235 4.155 ;
        RECT  3.225 3.685 4.865 4.155 ;
        RECT  2.760 3.455 3.225 4.155 ;
        RECT  0.545 3.685 2.760 4.155 ;
        RECT  0.165 3.115 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.360 2.360 5.445 2.700 ;
        RECT  5.130 1.245 5.360 3.225 ;
        RECT  3.285 1.245 5.130 1.475 ;
        RECT  1.520 2.995 5.130 3.225 ;
        RECT  1.905 0.495 4.610 0.725 ;
        RECT  2.935 0.955 3.285 1.475 ;
        RECT  1.675 0.495 1.905 1.440 ;
        RECT  0.465 1.210 1.675 1.440 ;
        RECT  0.235 0.635 0.465 1.440 ;
    END
END OA222D0BWP7T

MACRO OA222D1BWP7T
    CLASS CORE ;
    FOREIGN OA222D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 0.465 6.580 3.320 ;
        RECT  6.180 0.465 6.300 1.285 ;
        RECT  6.180 2.460 6.300 3.320 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.660 4.340 2.710 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.715 5.460 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.715 2.660 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.650 3.780 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.660 1.540 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.690 -0.235 6.720 0.235 ;
        RECT  5.460 -0.235 5.690 1.255 ;
        RECT  4.330 -0.235 5.460 0.235 ;
        RECT  3.950 -0.235 4.330 0.785 ;
        RECT  0.000 -0.235 3.950 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.770 3.685 6.720 4.155 ;
        RECT  5.390 2.850 5.770 4.155 ;
        RECT  3.370 3.685 5.390 4.155 ;
        RECT  3.140 2.840 3.370 4.155 ;
        RECT  0.570 3.685 3.140 4.155 ;
        RECT  0.340 2.940 0.570 4.155 ;
        RECT  0.000 3.685 0.340 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.700 1.660 5.930 2.620 ;
        RECT  5.045 2.380 5.700 2.620 ;
        RECT  4.805 2.380 5.045 3.170 ;
        RECT  4.740 0.465 4.970 1.275 ;
        RECT  3.830 2.940 4.805 3.170 ;
        RECT  2.445 1.015 4.740 1.275 ;
        RECT  3.600 2.380 3.830 3.170 ;
        RECT  2.625 2.380 3.600 2.610 ;
        RECT  2.010 0.480 3.505 0.765 ;
        RECT  2.300 2.380 2.625 3.170 ;
        RECT  1.030 2.940 2.300 3.170 ;
        RECT  1.780 0.480 2.010 1.290 ;
        RECT  0.570 0.480 1.780 0.765 ;
        RECT  1.030 1.020 1.345 1.250 ;
        RECT  0.800 1.020 1.030 3.170 ;
        RECT  0.340 0.480 0.570 1.290 ;
    END
END OA222D1BWP7T

MACRO OA222D2BWP7T
    CLASS CORE ;
    FOREIGN OA222D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 1.210 6.585 2.150 ;
        RECT  6.250 1.210 6.435 3.385 ;
        RECT  6.195 0.495 6.250 3.385 ;
        RECT  6.020 0.495 6.195 1.435 ;
        RECT  5.965 3.155 6.195 3.385 ;
        END
    END Z
    PIN C2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.715 4.340 2.150 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.715 5.460 2.150 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.660 2.150 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.715 3.220 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.660 1.540 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.040 -0.235 7.280 0.235 ;
        RECT  6.660 -0.235 7.040 0.895 ;
        RECT  5.610 -0.235 6.660 0.235 ;
        RECT  5.230 -0.235 5.610 1.200 ;
        RECT  4.180 -0.235 5.230 0.235 ;
        RECT  3.800 -0.235 4.180 0.785 ;
        RECT  0.000 -0.235 3.800 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.060 3.685 7.280 4.155 ;
        RECT  6.680 2.550 7.060 4.155 ;
        RECT  5.610 3.685 6.680 4.155 ;
        RECT  5.230 3.005 5.610 4.155 ;
        RECT  3.290 3.685 5.230 4.155 ;
        RECT  2.910 3.005 3.290 4.155 ;
        RECT  0.550 3.685 2.910 4.155 ;
        RECT  0.315 3.060 0.550 4.155 ;
        RECT  0.000 3.685 0.315 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.735 1.660 5.965 2.730 ;
        RECT  4.190 2.490 5.735 2.730 ;
        RECT  4.515 0.485 4.870 1.250 ;
        RECT  2.345 1.020 4.515 1.250 ;
        RECT  3.960 2.490 4.190 3.360 ;
        RECT  2.625 2.490 3.960 2.730 ;
        RECT  1.910 0.495 3.405 0.740 ;
        RECT  2.385 2.490 2.625 3.315 ;
        RECT  1.020 3.085 2.385 3.315 ;
        RECT  1.680 0.495 1.910 1.305 ;
        RECT  0.470 0.495 1.680 0.740 ;
        RECT  1.020 0.975 1.245 1.205 ;
        RECT  0.780 0.975 1.020 3.315 ;
        RECT  0.240 0.495 0.470 1.305 ;
    END
END OA222D2BWP7T

MACRO OA22D0BWP7T
    CLASS CORE ;
    FOREIGN OA22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.6030 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 0.845 4.340 3.400 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 2.280 0.450 2.710 ;
        RECT  0.140 1.770 0.420 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 2.330 3.285 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 1.820 3.270 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.820 1.590 2.100 ;
        RECT  1.310 1.695 1.540 2.100 ;
        RECT  0.650 1.820 1.310 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 -0.235 4.480 0.235 ;
        RECT  3.240 -0.235 3.580 1.130 ;
        RECT  0.520 -0.235 3.240 0.235 ;
        RECT  0.180 -0.235 0.520 1.130 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 3.685 4.480 4.155 ;
        RECT  2.960 3.455 3.300 4.155 ;
        RECT  0.520 3.685 2.960 4.155 ;
        RECT  0.180 3.075 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.535 1.360 3.765 3.215 ;
        RECT  2.025 1.360 3.535 1.590 ;
        RECT  1.460 2.985 3.535 3.215 ;
        RECT  2.750 0.900 2.860 1.130 ;
        RECT  2.520 0.465 2.750 1.130 ;
        RECT  1.205 0.465 2.520 0.695 ;
        RECT  1.795 0.925 2.025 1.590 ;
        RECT  0.975 0.465 1.205 1.185 ;
    END
END OA22D0BWP7T

MACRO OA22D1BWP7T
    CLASS CORE ;
    FOREIGN OA22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 0.495 4.905 3.300 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.340 1.660 1.570 2.150 ;
        RECT  0.700 1.770 1.340 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.660 3.780 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.715 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.175 -0.235 5.040 0.235 ;
        RECT  3.795 -0.235 4.175 0.740 ;
        RECT  1.265 -0.235 3.795 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.105 3.685 5.040 4.155 ;
        RECT  3.725 3.030 4.105 4.155 ;
        RECT  3.325 3.685 3.725 4.155 ;
        RECT  2.925 3.030 3.325 4.155 ;
        RECT  0.650 3.685 2.925 4.155 ;
        RECT  0.270 3.035 0.650 4.155 ;
        RECT  0.000 3.685 0.270 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.085 0.980 4.325 2.800 ;
        RECT  2.340 0.980 4.085 1.210 ;
        RECT  1.910 2.520 4.085 2.800 ;
        RECT  1.905 0.510 3.400 0.740 ;
        RECT  1.680 2.520 1.910 3.390 ;
        RECT  1.675 0.510 1.905 1.300 ;
        RECT  0.465 1.060 1.675 1.300 ;
        RECT  0.235 0.490 0.465 1.300 ;
    END
END OA22D1BWP7T

MACRO OA22D2BWP7T
    CLASS CORE ;
    FOREIGN OA22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 0.495 4.900 3.350 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.340 1.660 1.570 2.150 ;
        RECT  0.700 1.770 1.340 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.190 1.770 3.785 2.150 ;
        RECT  2.940 1.660 3.190 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.715 2.660 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.620 -0.235 6.160 0.235 ;
        RECT  5.240 -0.235 5.620 1.205 ;
        RECT  4.180 -0.235 5.240 0.235 ;
        RECT  3.800 -0.235 4.180 0.745 ;
        RECT  1.280 -0.235 3.800 0.235 ;
        RECT  0.900 -0.235 1.280 0.825 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.605 3.685 6.160 4.155 ;
        RECT  5.225 2.565 5.605 4.155 ;
        RECT  4.185 3.685 5.225 4.155 ;
        RECT  3.805 3.075 4.185 4.155 ;
        RECT  3.295 3.685 3.805 4.155 ;
        RECT  2.895 3.075 3.295 4.155 ;
        RECT  0.680 3.685 2.895 4.155 ;
        RECT  0.300 3.035 0.680 4.155 ;
        RECT  0.000 3.685 0.300 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.080 0.975 4.320 2.800 ;
        RECT  2.355 0.975 4.080 1.205 ;
        RECT  1.910 2.520 4.080 2.800 ;
        RECT  1.920 0.495 3.415 0.745 ;
        RECT  1.690 0.495 1.920 1.305 ;
        RECT  1.680 2.520 1.910 3.390 ;
        RECT  0.480 1.075 1.690 1.305 ;
        RECT  0.250 0.495 0.480 1.305 ;
    END
END OA22D2BWP7T

MACRO OA31D0BWP7T
    CLASS CORE ;
    FOREIGN OA31D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.875 4.340 3.355 ;
        RECT  3.950 0.875 4.060 1.105 ;
        RECT  3.950 3.125 4.060 3.355 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.770 2.150 2.210 ;
        RECT  1.820 1.770 2.100 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 1.540 2.710 ;
        RECT  1.240 2.360 1.260 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 1.010 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.560 -0.235 4.480 0.235 ;
        RECT  3.180 -0.235 3.560 1.075 ;
        RECT  0.000 -0.235 3.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 3.685 4.480 4.155 ;
        RECT  3.200 3.085 3.580 4.155 ;
        RECT  0.510 3.685 3.200 4.155 ;
        RECT  0.280 3.050 0.510 4.155 ;
        RECT  0.000 3.685 0.280 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.525 1.305 3.755 2.750 ;
        RECT  2.045 1.305 3.525 1.540 ;
        RECT  2.745 2.520 3.525 2.750 ;
        RECT  2.470 0.465 2.810 1.075 ;
        RECT  2.515 2.520 2.745 3.385 ;
        RECT  1.285 0.465 2.470 0.695 ;
        RECT  1.705 0.925 2.045 1.540 ;
        RECT  0.505 1.305 1.705 1.540 ;
        RECT  0.945 0.465 1.285 1.075 ;
        RECT  0.275 0.830 0.505 1.540 ;
    END
END OA31D0BWP7T

MACRO OA31D1BWP7T
    CLASS CORE ;
    FOREIGN OA31D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2129 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 0.545 4.340 2.620 ;
        RECT  4.060 0.545 4.245 3.390 ;
        RECT  3.905 0.545 4.060 0.775 ;
        RECT  4.015 2.375 4.060 3.390 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.650 3.225 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.670 2.145 2.100 ;
        RECT  1.820 1.670 2.100 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.680 1.540 2.710 ;
        RECT  1.210 1.680 1.255 2.035 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.675 0.980 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.485 -0.235 4.480 0.235 ;
        RECT  3.105 -0.235 3.485 0.790 ;
        RECT  0.000 -0.235 3.105 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.485 3.685 4.480 4.155 ;
        RECT  3.105 2.855 3.485 4.155 ;
        RECT  0.465 3.685 3.105 4.155 ;
        RECT  0.235 2.435 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.480 1.020 3.710 2.610 ;
        RECT  0.465 1.020 3.480 1.275 ;
        RECT  2.640 2.380 3.480 2.610 ;
        RECT  0.870 0.560 2.725 0.790 ;
        RECT  2.405 2.380 2.640 3.400 ;
        RECT  0.235 0.465 0.465 1.275 ;
    END
END OA31D1BWP7T

MACRO OA31D2BWP7T
    CLASS CORE ;
    FOREIGN OA31D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.3154 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.555 4.340 3.265 ;
        RECT  3.785 0.555 4.060 0.785 ;
        RECT  3.855 2.925 4.060 3.265 ;
        END
    END Z
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.670 3.225 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.670 2.100 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.730 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 -0.235 5.040 0.235 ;
        RECT  4.575 -0.235 4.805 1.265 ;
        RECT  3.420 -0.235 4.575 0.235 ;
        RECT  3.040 -0.235 3.420 0.770 ;
        RECT  0.000 -0.235 3.040 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 3.685 5.040 4.155 ;
        RECT  4.575 2.235 4.805 4.155 ;
        RECT  3.420 3.685 4.575 4.155 ;
        RECT  3.040 2.915 3.420 4.155 ;
        RECT  0.575 3.685 3.040 4.155 ;
        RECT  0.195 3.025 0.575 4.155 ;
        RECT  0.000 3.685 0.195 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.600 1.020 3.830 2.645 ;
        RECT  0.470 1.020 3.600 1.275 ;
        RECT  2.585 2.415 3.600 2.645 ;
        RECT  0.895 0.465 2.690 0.695 ;
        RECT  2.355 2.415 2.585 3.365 ;
        RECT  0.240 0.465 0.470 1.275 ;
    END
END OA31D2BWP7T

MACRO OA32D0BWP7T
    CLASS CORE ;
    FOREIGN OA32D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5520 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.015 5.460 3.330 ;
        RECT  5.040 1.015 5.180 1.245 ;
        RECT  4.660 3.100 5.180 3.330 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.770 3.220 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 4.340 2.160 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 2.230 2.100 3.270 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 1.770 1.540 3.270 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.765 -0.235 5.600 0.235 ;
        RECT  4.535 -0.235 4.765 0.540 ;
        RECT  0.000 -0.235 4.535 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.300 3.685 5.600 4.155 ;
        RECT  3.920 3.110 4.300 4.155 ;
        RECT  0.550 3.685 3.920 4.155 ;
        RECT  0.170 3.075 0.550 4.155 ;
        RECT  0.000 3.685 0.170 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.570 1.820 4.800 2.755 ;
        RECT  3.690 2.515 4.570 2.755 ;
        RECT  2.575 0.850 4.125 1.080 ;
        RECT  3.450 2.515 3.690 3.340 ;
        RECT  2.565 3.100 3.450 3.340 ;
        RECT  2.340 0.465 2.575 1.080 ;
        RECT  2.335 1.310 2.565 3.340 ;
        RECT  1.240 0.465 2.340 0.695 ;
        RECT  1.960 1.310 2.335 1.540 ;
        RECT  1.615 0.925 1.960 1.540 ;
        RECT  0.465 1.310 1.615 1.540 ;
        RECT  0.900 0.465 1.240 1.080 ;
        RECT  0.235 0.830 0.465 1.540 ;
    END
END OA32D0BWP7T

MACRO OA32D1BWP7T
    CLASS CORE ;
    FOREIGN OA32D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2198 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.130 0.495 5.460 2.750 ;
        RECT  4.945 2.470 5.130 2.750 ;
        RECT  4.715 2.470 4.945 3.280 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.660 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.660 3.810 2.710 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.680 2.150 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.680 1.545 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.615 -0.235 5.600 0.235 ;
        RECT  4.365 -0.235 4.615 0.555 ;
        RECT  3.405 -0.235 4.365 0.235 ;
        RECT  3.060 -0.235 3.405 0.770 ;
        RECT  0.000 -0.235 3.060 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.195 3.685 5.600 4.155 ;
        RECT  3.835 3.415 4.195 4.155 ;
        RECT  0.465 3.685 3.835 4.155 ;
        RECT  0.235 3.020 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.360 1.725 4.760 1.955 ;
        RECT  4.130 1.725 4.360 3.180 ;
        RECT  2.625 1.015 4.130 1.275 ;
        RECT  2.615 2.950 4.130 3.180 ;
        RECT  2.395 0.465 2.625 1.275 ;
        RECT  2.380 2.950 2.615 3.320 ;
        RECT  1.185 0.465 2.395 0.695 ;
        RECT  1.000 3.090 2.380 3.320 ;
        RECT  1.615 0.925 1.960 1.310 ;
        RECT  1.000 1.070 1.615 1.310 ;
        RECT  0.955 0.465 1.185 0.840 ;
        RECT  0.755 1.070 1.000 3.320 ;
        RECT  0.465 1.070 0.755 1.310 ;
        RECT  0.235 0.495 0.465 1.310 ;
    END
END OA32D1BWP7T

MACRO OA32D2BWP7T
    CLASS CORE ;
    FOREIGN OA32D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.775 1.165 6.020 2.750 ;
        RECT  5.765 0.495 5.775 2.750 ;
        RECT  5.740 0.495 5.765 3.280 ;
        RECT  5.530 0.495 5.740 1.470 ;
        RECT  5.535 2.415 5.740 3.280 ;
        END
    END Z
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.660 3.220 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.660 3.810 2.710 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.680 2.150 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.680 1.545 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.505 -0.235 6.720 0.235 ;
        RECT  6.255 -0.235 6.505 1.240 ;
        RECT  5.055 -0.235 6.255 0.235 ;
        RECT  4.805 -0.235 5.055 1.240 ;
        RECT  3.405 -0.235 4.805 0.235 ;
        RECT  3.060 -0.235 3.405 0.770 ;
        RECT  0.000 -0.235 3.060 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 3.685 6.720 4.155 ;
        RECT  6.250 2.440 6.490 4.155 ;
        RECT  5.050 3.685 6.250 4.155 ;
        RECT  4.810 2.440 5.050 4.155 ;
        RECT  4.195 3.685 4.810 4.155 ;
        RECT  3.835 3.415 4.195 4.155 ;
        RECT  0.465 3.685 3.835 4.155 ;
        RECT  0.235 3.020 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.495 1.670 5.290 1.900 ;
        RECT  4.265 1.670 4.495 3.180 ;
        RECT  2.615 2.950 4.265 3.180 ;
        RECT  3.835 0.465 4.065 1.275 ;
        RECT  2.625 1.015 3.835 1.275 ;
        RECT  2.395 0.465 2.625 1.275 ;
        RECT  2.380 2.950 2.615 3.320 ;
        RECT  1.185 0.465 2.395 0.695 ;
        RECT  1.000 3.090 2.380 3.320 ;
        RECT  1.615 0.925 1.960 1.310 ;
        RECT  1.000 1.070 1.615 1.310 ;
        RECT  0.955 0.465 1.185 0.840 ;
        RECT  0.755 1.070 1.000 3.320 ;
        RECT  0.465 1.070 0.755 1.310 ;
        RECT  0.235 0.495 0.465 1.310 ;
    END
END OA32D2BWP7T

MACRO OA33D0BWP7T
    CLASS CORE ;
    FOREIGN OA33D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 0.780 5.460 3.320 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 1.770 3.780 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.770 4.340 2.725 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.770 2.150 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.770 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.650 -0.235 5.600 0.235 ;
        RECT  4.310 -0.235 4.650 0.465 ;
        RECT  3.460 -0.235 4.310 0.235 ;
        RECT  3.120 -0.235 3.460 0.465 ;
        RECT  0.000 -0.235 3.120 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 3.685 5.600 4.155 ;
        RECT  4.180 3.455 4.540 4.155 ;
        RECT  0.545 3.685 4.180 4.155 ;
        RECT  0.165 3.155 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.620 1.635 4.900 3.225 ;
        RECT  3.080 2.985 4.620 3.225 ;
        RECT  2.645 1.095 4.035 1.335 ;
        RECT  2.840 2.985 3.080 3.325 ;
        RECT  1.020 3.095 2.840 3.325 ;
        RECT  2.415 0.465 2.645 1.335 ;
        RECT  1.260 0.465 2.415 0.695 ;
        RECT  1.640 0.930 1.980 1.540 ;
        RECT  1.020 1.310 1.640 1.540 ;
        RECT  0.920 0.465 1.260 1.080 ;
        RECT  0.780 1.310 1.020 3.325 ;
        RECT  0.535 1.310 0.780 1.540 ;
        RECT  0.195 0.905 0.535 1.540 ;
    END
END OA33D0BWP7T

MACRO OA33D1BWP7T
    CLASS CORE ;
    FOREIGN OA33D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2472 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 1.170 6.020 2.680 ;
        RECT  5.740 0.495 5.760 2.680 ;
        RECT  5.530 0.495 5.740 1.440 ;
        RECT  5.540 2.440 5.740 2.680 ;
        RECT  5.310 2.440 5.540 3.435 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 1.210 3.220 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.825 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.725 4.615 1.955 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.680 2.100 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.735 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.465 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.040 -0.235 6.160 0.235 ;
        RECT  4.810 -0.235 5.040 1.260 ;
        RECT  3.525 -0.235 4.810 0.235 ;
        RECT  3.150 -0.235 3.525 0.465 ;
        RECT  0.000 -0.235 3.150 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.885 3.685 6.160 4.155 ;
        RECT  4.505 2.945 4.885 4.155 ;
        RECT  0.560 3.685 4.505 4.155 ;
        RECT  0.180 3.025 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.080 1.735 5.335 1.965 ;
        RECT  4.850 1.735 5.080 2.670 ;
        RECT  2.585 2.430 4.850 2.670 ;
        RECT  2.625 0.695 4.410 0.935 ;
        RECT  2.395 0.465 2.625 0.935 ;
        RECT  2.355 1.190 2.585 3.415 ;
        RECT  1.245 0.465 2.395 0.705 ;
        RECT  1.965 1.190 2.355 1.430 ;
        RECT  1.610 0.935 1.965 1.430 ;
        RECT  0.465 1.190 1.610 1.430 ;
        RECT  0.890 0.465 1.245 0.840 ;
        RECT  0.235 0.495 0.465 1.430 ;
    END
END OA33D1BWP7T

MACRO OA33D2BWP7T
    CLASS CORE ;
    FOREIGN OA33D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.3072 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 1.170 6.020 2.485 ;
        RECT  5.740 0.495 5.760 2.485 ;
        RECT  5.530 0.495 5.740 1.440 ;
        RECT  5.540 2.245 5.740 2.485 ;
        RECT  5.310 2.245 5.540 3.405 ;
        END
    END Z
    PIN B3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 1.210 3.220 2.150 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.825 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.725 4.615 1.955 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.680 2.100 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.735 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.465 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.560 -0.235 6.720 0.235 ;
        RECT  6.175 -0.235 6.560 0.935 ;
        RECT  5.040 -0.235 6.175 0.235 ;
        RECT  4.810 -0.235 5.040 1.260 ;
        RECT  3.525 -0.235 4.810 0.235 ;
        RECT  3.150 -0.235 3.525 0.465 ;
        RECT  0.000 -0.235 3.150 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.345 3.685 6.720 4.155 ;
        RECT  5.965 2.750 6.345 4.155 ;
        RECT  4.885 3.685 5.965 4.155 ;
        RECT  4.505 2.945 4.885 4.155 ;
        RECT  0.560 3.685 4.505 4.155 ;
        RECT  0.180 3.025 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.080 1.670 5.335 1.900 ;
        RECT  4.850 1.670 5.080 2.670 ;
        RECT  2.585 2.430 4.850 2.670 ;
        RECT  2.625 0.695 4.410 0.935 ;
        RECT  2.395 0.465 2.625 0.935 ;
        RECT  2.355 1.190 2.585 3.415 ;
        RECT  1.245 0.465 2.395 0.705 ;
        RECT  1.965 1.190 2.355 1.430 ;
        RECT  1.610 0.935 1.965 1.430 ;
        RECT  0.465 1.190 1.610 1.430 ;
        RECT  0.890 0.465 1.245 0.840 ;
        RECT  0.235 0.495 0.465 1.430 ;
    END
END OA33D2BWP7T

MACRO OAI211D0BWP7T
    CLASS CORE ;
    FOREIGN OAI211D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9787 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 2.380 3.125 3.345 ;
        RECT  2.660 2.380 2.895 2.660 ;
        RECT  2.380 0.775 2.660 2.660 ;
        RECT  2.120 0.775 2.380 1.005 ;
        RECT  1.185 2.380 2.380 2.660 ;
        RECT  0.955 2.380 1.185 3.345 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.465 2.710 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.540 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.210 3.220 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.260 2.150 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 -0.235 3.360 0.235 ;
        RECT  0.160 -0.235 0.540 1.045 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 3.685 3.360 4.155 ;
        RECT  1.605 3.045 1.985 4.155 ;
        RECT  0.550 3.685 1.605 4.155 ;
        RECT  0.170 3.045 0.550 4.155 ;
        RECT  0.000 3.685 0.170 4.155 ;
        END
    END VDD
END OAI211D0BWP7T

MACRO OAI211D1BWP7T
    CLASS CORE ;
    FOREIGN OAI211D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.9374 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 2.425 3.125 3.235 ;
        RECT  2.660 2.425 2.895 2.655 ;
        RECT  2.380 0.960 2.660 2.655 ;
        RECT  0.960 0.960 2.380 1.190 ;
        RECT  0.960 2.940 1.240 3.170 ;
        RECT  0.730 0.960 0.960 3.170 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.215 1.610 1.540 2.710 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.210 3.220 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.610 2.115 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 -0.235 3.360 0.235 ;
        RECT  0.155 -0.235 0.535 0.835 ;
        RECT  0.000 -0.235 0.155 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 3.685 3.360 4.155 ;
        RECT  1.605 2.940 1.985 4.155 ;
        RECT  0.465 3.685 1.605 4.155 ;
        RECT  0.235 2.685 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.400 0.500 3.180 0.730 ;
    END
END OAI211D1BWP7T

MACRO OAI211D2BWP7T
    CLASS CORE ;
    FOREIGN OAI211D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.2994 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 0.925 6.020 3.120 ;
        RECT  3.480 0.925 5.740 1.155 ;
        RECT  4.205 2.890 5.740 3.120 ;
        RECT  3.930 2.790 4.205 3.120 ;
        RECT  0.895 2.790 3.930 3.020 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 1.770 2.100 2.150 ;
        END
    END C
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 1.260 2.805 1.870 ;
        RECT  0.700 1.260 2.575 1.540 ;
        RECT  0.470 1.260 0.700 1.995 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 1.680 4.950 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.685 5.495 2.560 ;
        RECT  3.780 2.330 5.180 2.560 ;
        RECT  3.500 1.665 3.780 2.560 ;
        RECT  3.290 1.665 3.500 1.895 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.780 -0.235 6.160 0.235 ;
        RECT  1.440 -0.235 1.780 0.565 ;
        RECT  0.000 -0.235 1.440 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 3.685 6.160 4.155 ;
        RECT  5.640 3.350 5.980 4.155 ;
        RECT  3.420 3.685 5.640 4.155 ;
        RECT  3.080 3.250 3.420 4.155 ;
        RECT  1.990 3.685 3.080 4.155 ;
        RECT  1.610 3.250 1.990 4.155 ;
        RECT  0.520 3.685 1.610 4.155 ;
        RECT  0.180 2.310 0.520 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.045 0.465 5.980 0.695 ;
        RECT  2.815 0.465 3.045 1.030 ;
        RECT  0.180 0.800 2.815 1.030 ;
    END
END OAI211D2BWP7T

MACRO OAI21D0BWP7T
    CLASS CORE ;
    FOREIGN OAI21D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.6433 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 3.015 1.875 3.245 ;
        RECT  0.980 0.980 1.240 1.210 ;
        RECT  0.700 0.980 0.980 3.245 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2070 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.350 1.210 2.660 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.770 2.100 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 -0.235 2.800 0.235 ;
        RECT  2.330 -0.235 2.570 0.585 ;
        RECT  0.000 -0.235 2.330 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.620 3.685 2.800 4.155 ;
        RECT  2.240 3.020 2.620 4.155 ;
        RECT  0.465 3.685 2.240 4.155 ;
        RECT  0.235 2.955 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.675 0.505 1.905 1.280 ;
        RECT  0.465 0.505 1.675 0.735 ;
        RECT  0.235 0.505 0.465 1.265 ;
    END
END OAI21D0BWP7T

MACRO OAI21D1BWP7T
    CLASS CORE ;
    FOREIGN OAI21D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.8552 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.535 2.380 2.765 3.345 ;
        RECT  0.980 2.380 2.535 2.660 ;
        RECT  1.095 0.925 1.325 1.770 ;
        RECT  0.980 1.540 1.095 1.770 ;
        RECT  0.700 1.540 0.980 3.190 ;
        RECT  0.320 2.960 0.700 3.190 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.720 3.220 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.100 2.150 ;
        RECT  1.570 1.730 1.820 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.690 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 -0.235 3.360 0.235 ;
        RECT  2.535 -0.235 2.770 1.265 ;
        RECT  0.000 -0.235 2.535 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 3.685 3.360 4.155 ;
        RECT  1.815 2.925 2.045 4.155 ;
        RECT  0.000 3.685 1.815 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.815 0.465 2.045 0.910 ;
        RECT  0.605 0.465 1.815 0.695 ;
        RECT  0.375 0.465 0.605 1.275 ;
    END
END OAI21D1BWP7T

MACRO OAI21D2BWP7T
    CLASS CORE ;
    FOREIGN OAI21D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.5665 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 0.940 4.900 3.120 ;
        RECT  2.350 0.940 4.620 1.170 ;
        RECT  0.905 2.890 4.620 3.120 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.735 1.540 2.150 ;
        END
    END B
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.135 1.590 4.365 2.660 ;
        RECT  2.405 2.380 4.135 2.660 ;
        RECT  2.170 1.700 2.405 2.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 1.780 3.830 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 -0.235 5.040 0.235 ;
        RECT  0.905 -0.235 1.245 0.670 ;
        RECT  0.000 -0.235 0.905 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.880 3.685 5.040 4.155 ;
        RECT  4.500 3.360 4.880 4.155 ;
        RECT  2.035 3.685 4.500 4.155 ;
        RECT  1.630 3.350 2.035 4.155 ;
        RECT  0.465 3.685 1.630 4.155 ;
        RECT  0.235 2.210 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.925 0.465 4.890 0.695 ;
        RECT  1.695 0.465 1.925 1.130 ;
        RECT  0.180 0.900 1.695 1.130 ;
    END
END OAI21D2BWP7T

MACRO OAI221D0BWP7T
    CLASS CORE ;
    FOREIGN OAI221D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9858 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 2.940 3.835 3.220 ;
        RECT  1.540 0.955 2.900 1.185 ;
        RECT  1.310 0.955 1.540 3.220 ;
        RECT  0.945 2.940 1.310 3.220 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 0.985 0.450 2.150 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 1.705 1.080 2.045 ;
        RECT  0.700 1.705 0.980 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.030 1.910 4.265 2.660 ;
        RECT  1.845 2.380 4.030 2.660 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.720 2.695 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 3.780 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.560 -0.235 4.480 0.235 ;
        RECT  0.180 -0.235 0.560 0.690 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.505 3.685 4.480 4.155 ;
        RECT  2.135 3.455 2.505 4.155 ;
        RECT  0.560 3.685 2.135 4.155 ;
        RECT  0.180 3.120 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.010 0.480 4.240 1.240 ;
        RECT  0.905 0.480 4.010 0.710 ;
    END
END OAI221D0BWP7T

MACRO OAI221D1BWP7T
    CLASS CORE ;
    FOREIGN OAI221D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.9374 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 1.015 4.900 3.315 ;
        RECT  3.800 1.015 4.575 1.245 ;
        RECT  3.830 3.085 4.575 3.315 ;
        RECT  3.600 2.440 3.830 3.315 ;
        RECT  1.190 2.440 3.600 2.670 ;
        RECT  0.960 2.440 1.190 3.350 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.705 0.450 2.710 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.670 1.540 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.665 2.660 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.725 4.345 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 -0.235 5.040 0.235 ;
        RECT  0.240 -0.235 0.470 1.205 ;
        RECT  0.000 -0.235 0.240 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.370 3.685 5.040 4.155 ;
        RECT  3.130 3.000 3.370 4.155 ;
        RECT  2.395 3.685 3.130 4.155 ;
        RECT  2.155 3.000 2.395 4.155 ;
        RECT  0.550 3.685 2.155 4.155 ;
        RECT  0.170 3.040 0.550 4.155 ;
        RECT  0.000 3.685 0.170 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.365 0.535 4.860 0.765 ;
        RECT  3.135 0.535 3.365 1.245 ;
        RECT  1.625 1.015 3.135 1.245 ;
        RECT  1.245 0.535 2.685 0.765 ;
        RECT  0.905 0.535 1.245 1.235 ;
    END
END OAI221D1BWP7T

MACRO OAI221D2BWP7T
    CLASS CORE ;
    FOREIGN OAI221D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 5.0472 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.460 0.925 8.660 1.155 ;
        RECT  5.460 2.940 8.550 3.220 ;
        RECT  5.180 0.925 5.460 3.220 ;
        RECT  4.825 2.940 5.180 3.220 ;
        RECT  4.595 2.445 4.825 3.220 ;
        RECT  1.985 2.940 4.595 3.220 ;
        RECT  1.755 2.380 1.985 3.220 ;
        RECT  0.465 2.380 1.755 2.610 ;
        RECT  0.235 2.380 0.465 3.410 ;
        END
    END ZN
    PIN C
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.540 2.150 ;
        END
    END C
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.635 4.665 1.865 ;
        RECT  4.060 1.635 4.340 2.660 ;
        RECT  2.660 2.380 4.060 2.660 ;
        RECT  2.380 1.665 2.660 2.660 ;
        RECT  1.970 1.665 2.380 1.895 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.590 3.780 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.655 7.700 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.030 1.580 8.265 2.660 ;
        RECT  5.985 2.380 8.030 2.660 ;
        RECT  5.755 1.580 5.985 2.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 -0.235 8.960 0.235 ;
        RECT  0.930 -0.235 1.280 0.670 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.200 3.685 8.960 4.155 ;
        RECT  6.800 3.455 7.200 4.155 ;
        RECT  3.540 3.685 6.800 4.155 ;
        RECT  3.160 3.455 3.540 4.155 ;
        RECT  1.230 3.685 3.160 4.155 ;
        RECT  1.000 2.900 1.230 4.155 ;
        RECT  0.000 3.685 1.000 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.420 0.465 7.900 0.695 ;
        RECT  0.180 0.925 4.920 1.155 ;
    END
END OAI221D2BWP7T

MACRO OAI222D0BWP7T
    CLASS CORE ;
    FOREIGN OAI222D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9756 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 2.970 4.360 3.200 ;
        RECT  3.180 0.990 3.520 1.385 ;
        RECT  0.980 1.155 3.180 1.385 ;
        RECT  0.700 1.155 0.980 3.200 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.615 1.540 2.710 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.795 1.770 2.100 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 1.740 4.805 2.660 ;
        RECT  2.750 2.380 4.575 2.660 ;
        RECT  2.410 2.335 2.750 2.660 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 1.665 3.270 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 4.340 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 -0.235 5.040 0.235 ;
        RECT  0.945 -0.235 1.325 0.465 ;
        RECT  0.000 -0.235 0.945 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.105 3.685 5.040 4.155 ;
        RECT  2.750 3.430 3.105 4.155 ;
        RECT  0.465 3.685 2.750 4.155 ;
        RECT  0.230 2.965 0.465 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.575 0.465 4.805 1.275 ;
        RECT  2.085 0.465 4.575 0.705 ;
        RECT  1.855 0.465 2.085 0.925 ;
        RECT  0.465 0.695 1.855 0.925 ;
        RECT  0.235 0.695 0.465 1.260 ;
    END
END OAI222D0BWP7T

MACRO OAI222D1BWP7T
    CLASS CORE ;
    FOREIGN OAI222D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.0110 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 2.380 5.365 3.420 ;
        RECT  4.900 2.380 5.135 2.660 ;
        RECT  4.620 0.925 4.900 2.660 ;
        RECT  4.415 0.925 4.620 1.265 ;
        RECT  2.870 2.380 4.620 2.660 ;
        RECT  2.640 2.380 2.870 3.235 ;
        RECT  1.600 3.005 2.640 3.235 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.540 2.150 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.725 0.455 2.710 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.725 2.100 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4050 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.740 3.220 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4050 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.745 4.340 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4131 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.210 5.460 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.295 -0.235 5.600 0.235 ;
        RECT  0.835 -0.235 1.295 0.780 ;
        RECT  0.000 -0.235 0.835 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.815 3.685 5.600 4.155 ;
        RECT  3.435 2.890 3.815 4.155 ;
        RECT  0.545 3.685 3.435 4.155 ;
        RECT  0.160 3.010 0.545 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.040 0.465 5.425 0.695 ;
        RECT  3.800 0.465 4.040 1.370 ;
        RECT  2.685 1.140 3.800 1.370 ;
        RECT  1.905 0.465 3.440 0.695 ;
        RECT  2.340 0.960 2.685 1.370 ;
        RECT  1.675 0.465 1.905 1.275 ;
        RECT  0.465 1.045 1.675 1.275 ;
        RECT  0.235 0.465 0.465 1.275 ;
    END
END OAI222D1BWP7T

MACRO OAI222D2BWP7T
    CLASS CORE ;
    FOREIGN OAI222D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.7294 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.805 1.015 9.940 3.020 ;
        RECT  9.660 0.490 9.805 3.020 ;
        RECT  9.575 0.490 9.660 1.245 ;
        RECT  1.575 2.790 9.660 3.020 ;
        RECT  6.640 1.015 9.575 1.245 ;
        END
    END ZN
    PIN C2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 1.675 2.195 2.100 ;
        END
    END C2
    PIN C1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.655 1.675 2.885 2.560 ;
        RECT  0.450 2.330 2.655 2.560 ;
        RECT  0.420 1.630 0.450 2.560 ;
        RECT  0.140 1.630 0.420 2.710 ;
        END
    END C1
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 1.695 5.070 2.100 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.595 6.020 2.560 ;
        RECT  3.780 2.330 5.740 2.560 ;
        RECT  3.475 1.645 3.780 2.560 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.100 1.575 9.380 2.560 ;
        RECT  7.140 2.330 9.100 2.560 ;
        RECT  6.860 1.625 7.140 2.560 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.845 1.675 8.870 2.100 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.700 -0.235 10.080 0.235 ;
        RECT  2.320 -0.235 2.700 0.765 ;
        RECT  1.255 -0.235 2.320 0.235 ;
        RECT  0.875 -0.235 1.255 0.765 ;
        RECT  0.000 -0.235 0.875 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.670 3.685 10.080 4.155 ;
        RECT  9.315 3.250 9.670 4.155 ;
        RECT  7.040 3.685 9.315 4.155 ;
        RECT  6.580 3.250 7.040 4.155 ;
        RECT  6.140 3.685 6.580 4.155 ;
        RECT  5.800 3.250 6.140 4.155 ;
        RECT  3.280 3.685 5.800 4.155 ;
        RECT  2.885 3.250 3.280 4.155 ;
        RECT  0.540 3.685 2.885 4.155 ;
        RECT  0.160 3.010 0.540 4.155 ;
        RECT  0.000 3.685 0.160 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.780 0.535 9.140 0.765 ;
        RECT  3.345 1.015 6.280 1.245 ;
        RECT  3.115 0.490 3.345 1.245 ;
        RECT  1.905 1.015 3.115 1.245 ;
        RECT  1.675 0.490 1.905 1.245 ;
        RECT  0.520 1.015 1.675 1.245 ;
        RECT  0.180 0.535 0.520 1.245 ;
    END
END OAI222D2BWP7T

MACRO OAI22D0BWP7T
    CLASS CORE ;
    FOREIGN OAI22D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.7871 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.870 2.100 2.995 ;
        RECT  1.505 0.870 1.820 1.100 ;
        RECT  1.610 2.765 1.820 2.995 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.455 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 0.985 3.220 2.660 ;
        RECT  2.665 2.380 2.910 2.660 ;
        RECT  2.435 2.380 2.665 3.455 ;
        RECT  1.380 3.225 2.435 3.455 ;
        RECT  1.150 2.410 1.380 3.455 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.375 1.210 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.590 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.190 -0.235 3.360 0.235 ;
        RECT  2.810 -0.235 3.190 0.710 ;
        RECT  0.535 -0.235 2.810 0.235 ;
        RECT  0.155 -0.235 0.535 0.845 ;
        RECT  0.000 -0.235 0.155 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 3.685 3.360 4.155 ;
        RECT  2.895 3.020 3.125 4.155 ;
        RECT  0.560 3.685 2.895 4.155 ;
        RECT  0.180 3.115 0.560 4.155 ;
        RECT  0.000 3.685 0.180 4.155 ;
        END
    END VDD
END OAI22D0BWP7T

MACRO OAI22D1BWP7T
    CLASS CORE ;
    FOREIGN OAI22D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.1026 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 0.965 3.685 3.220 ;
        RECT  2.590 0.965 3.455 1.195 ;
        RECT  0.200 2.940 3.455 3.220 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.655 1.540 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.630 0.465 2.710 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.745 2.660 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.630 3.220 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.235 3.920 0.235 ;
        RECT  0.940 -0.235 1.310 0.775 ;
        RECT  0.000 -0.235 0.940 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.185 3.685 3.920 4.155 ;
        RECT  1.845 3.455 2.185 4.155 ;
        RECT  0.000 3.685 1.845 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.005 0.505 3.755 0.735 ;
        RECT  1.775 0.505 2.005 1.275 ;
        RECT  0.485 1.045 1.775 1.275 ;
        RECT  0.255 0.465 0.485 1.275 ;
    END
END OAI22D1BWP7T

MACRO OAI22D2BWP7T
    CLASS CORE ;
    FOREIGN OAI22D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.6344 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 0.995 6.580 3.070 ;
        RECT  3.980 0.995 6.300 1.225 ;
        RECT  1.680 2.840 6.300 3.070 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.570 3.220 2.610 ;
        RECT  0.980 2.380 2.855 2.610 ;
        RECT  0.700 1.570 0.980 2.610 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.575 2.250 2.150 ;
        END
    END B1
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.570 6.020 2.610 ;
        RECT  3.780 2.380 5.740 2.610 ;
        RECT  3.500 1.570 3.780 2.610 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.415 1.575 5.460 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 -0.235 6.720 0.235 ;
        RECT  2.420 -0.235 2.820 0.670 ;
        RECT  1.305 -0.235 2.420 0.235 ;
        RECT  0.905 -0.235 1.305 0.670 ;
        RECT  0.000 -0.235 0.905 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 3.685 6.720 4.155 ;
        RECT  5.990 3.300 6.335 4.155 ;
        RECT  3.515 3.685 5.990 4.155 ;
        RECT  3.145 3.300 3.515 4.155 ;
        RECT  0.470 3.685 3.145 4.155 ;
        RECT  0.240 2.475 0.470 4.155 ;
        RECT  0.000 3.685 0.240 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.505 0.535 6.480 0.765 ;
        RECT  3.275 0.535 3.505 1.275 ;
        RECT  1.965 1.035 3.275 1.275 ;
        RECT  1.735 0.465 1.965 1.275 ;
        RECT  0.470 1.035 1.735 1.275 ;
        RECT  0.240 0.465 0.470 1.275 ;
    END
END OAI22D2BWP7T

MACRO OAI31D0BWP7T
    CLASS CORE ;
    FOREIGN OAI31D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.9098 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.980 2.660 3.245 ;
        RECT  0.180 0.980 2.380 1.210 ;
        RECT  2.085 3.015 2.380 3.245 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.900 1.770 3.220 2.710 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.770 2.105 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.765 1.540 2.225 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.465 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.235 3.360 0.235 ;
        RECT  2.895 -0.235 3.125 1.245 ;
        RECT  0.000 -0.235 2.895 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 3.685 3.360 4.155 ;
        RECT  2.895 3.035 3.125 4.155 ;
        RECT  0.545 3.685 2.895 4.155 ;
        RECT  0.165 3.085 0.545 4.155 ;
        RECT  0.000 3.685 0.165 4.155 ;
        END
    END VDD
END OAI31D0BWP7T

MACRO OAI31D1BWP7T
    CLASS CORE ;
    FOREIGN OAI31D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.9831 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 3.040 2.780 3.270 ;
        RECT  1.820 1.020 2.100 3.270 ;
        RECT  0.525 1.020 1.820 1.275 ;
        RECT  0.295 0.465 0.525 1.275 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 3.780 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 1.630 2.660 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.755 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.630 0.465 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 -0.235 3.920 0.235 ;
        RECT  3.260 -0.235 3.495 1.290 ;
        RECT  0.000 -0.235 3.260 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 3.685 3.920 4.155 ;
        RECT  3.265 2.435 3.495 4.155 ;
        RECT  0.600 3.685 3.265 4.155 ;
        RECT  0.220 3.020 0.600 4.155 ;
        RECT  0.000 3.685 0.220 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.515 0.465 2.745 1.275 ;
        RECT  0.950 0.465 2.515 0.725 ;
    END
END OAI31D1BWP7T

MACRO OAI31D2BWP7T
    CLASS CORE ;
    FOREIGN OAI31D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.9511 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 0.925 5.655 1.155 ;
        RECT  2.630 3.225 4.235 3.455 ;
        RECT  2.400 2.940 2.630 3.455 ;
        RECT  1.540 2.940 2.400 3.225 ;
        RECT  1.915 0.925 2.145 1.515 ;
        RECT  1.540 1.285 1.915 1.515 ;
        RECT  1.260 1.285 1.540 3.225 ;
        RECT  0.955 2.885 1.260 3.225 ;
        END
    END ZN
    PIN B
        ANTENNAGATEAREA 0.8280 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.730 1.000 2.150 ;
        END
    END B
    PIN A3
        ANTENNAGATEAREA 0.8046 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.290 2.380 6.070 2.660 ;
        RECT  4.985 2.305 5.290 2.660 ;
        RECT  4.200 2.305 4.985 2.535 ;
        RECT  3.860 1.845 4.200 2.535 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 1.490 6.580 3.220 ;
        RECT  6.205 1.490 6.300 1.720 ;
        RECT  4.770 2.940 6.300 3.220 ;
        RECT  4.540 2.765 4.770 3.220 ;
        RECT  3.220 2.765 4.540 2.995 ;
        RECT  2.940 1.845 3.220 2.995 ;
        RECT  2.835 1.845 2.940 2.185 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8064 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.540 1.385 5.880 2.130 ;
        RECT  2.605 1.385 5.540 1.615 ;
        RECT  2.375 1.385 2.605 2.000 ;
        RECT  2.100 1.770 2.375 2.000 ;
        RECT  1.820 1.770 2.100 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 -0.235 6.720 0.235 ;
        RECT  0.995 -0.235 1.225 0.520 ;
        RECT  0.000 -0.235 0.995 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.540 3.685 6.720 4.155 ;
        RECT  6.200 3.455 6.540 4.155 ;
        RECT  2.025 3.685 6.200 4.155 ;
        RECT  1.645 3.455 2.025 4.155 ;
        RECT  0.465 3.685 1.645 4.155 ;
        RECT  0.235 2.435 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.685 0.465 6.390 0.695 ;
        RECT  1.455 0.465 1.685 0.985 ;
        RECT  0.175 0.750 1.455 0.985 ;
    END
END OAI31D2BWP7T

MACRO OAI32D0BWP7T
    CLASS CORE ;
    FOREIGN OAI32D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.790 2.660 3.370 ;
        RECT  2.010 1.790 2.380 2.100 ;
        RECT  1.770 0.925 2.010 2.100 ;
        RECT  1.670 0.925 1.770 1.540 ;
        RECT  0.510 1.310 1.670 1.540 ;
        RECT  0.280 0.830 0.510 1.540 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.770 3.220 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 4.340 2.185 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 2.330 2.145 3.270 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 2.330 1.540 3.270 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.980 2.220 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.485 -0.235 4.480 0.235 ;
        RECT  3.105 -0.235 3.485 1.075 ;
        RECT  0.000 -0.235 3.105 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.210 3.685 4.480 4.155 ;
        RECT  3.830 3.135 4.210 4.155 ;
        RECT  0.585 3.685 3.830 4.155 ;
        RECT  0.205 3.085 0.585 4.155 ;
        RECT  0.000 3.685 0.205 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.900 0.825 4.130 1.540 ;
        RECT  2.690 1.310 3.900 1.540 ;
        RECT  2.460 0.465 2.690 1.540 ;
        RECT  1.290 0.465 2.460 0.695 ;
        RECT  0.950 0.465 1.290 1.080 ;
    END
END OAI32D0BWP7T

MACRO OAI32D1BWP7T
    CLASS CORE ;
    FOREIGN OAI32D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.2680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 2.410 2.705 3.270 ;
        RECT  0.985 3.040 2.475 3.270 ;
        RECT  1.675 0.925 2.030 1.380 ;
        RECT  0.985 1.150 1.675 1.380 ;
        RECT  0.755 1.150 0.985 3.270 ;
        RECT  0.700 1.150 0.755 2.835 ;
        RECT  0.500 1.150 0.700 1.380 ;
        RECT  0.270 0.480 0.500 1.380 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.635 3.220 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.690 4.340 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.655 2.660 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.610 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.610 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 -0.235 4.480 0.235 ;
        RECT  3.120 -0.235 3.500 0.855 ;
        RECT  0.000 -0.235 3.120 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 3.685 4.480 4.155 ;
        RECT  3.910 2.500 4.140 4.155 ;
        RECT  0.500 3.685 3.910 4.155 ;
        RECT  0.270 2.995 0.500 4.155 ;
        RECT  0.000 3.685 0.270 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.910 0.495 4.140 1.400 ;
        RECT  2.700 1.170 3.910 1.400 ;
        RECT  2.470 0.465 2.700 1.400 ;
        RECT  1.300 0.465 2.470 0.695 ;
        RECT  0.960 0.465 1.300 0.870 ;
    END
END OAI32D1BWP7T

MACRO OAI32D2BWP7T
    CLASS CORE ;
    FOREIGN OAI32D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.400 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.0996 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 0.955 8.260 2.855 ;
        RECT  3.825 0.955 7.980 1.185 ;
        RECT  7.125 2.605 7.980 2.855 ;
        RECT  3.585 0.955 3.825 2.535 ;
        RECT  3.335 2.305 3.585 2.535 ;
        RECT  3.105 2.305 3.335 3.070 ;
        RECT  1.510 2.840 3.105 3.070 ;
        END
    END ZN
    PIN B2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.740 2.110 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.645 1.690 2.875 2.610 ;
        RECT  0.980 2.380 2.645 2.610 ;
        RECT  0.700 1.700 0.980 2.610 ;
        RECT  0.140 1.700 0.700 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.605 7.700 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.655 6.020 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.8532 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.675 4.900 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.705 -0.235 8.400 0.235 ;
        RECT  2.325 -0.235 2.705 0.885 ;
        RECT  1.265 -0.235 2.325 0.235 ;
        RECT  0.885 -0.235 1.265 0.880 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.625 3.685 8.400 4.155 ;
        RECT  4.285 3.225 4.625 4.155 ;
        RECT  3.150 3.685 4.285 4.155 ;
        RECT  2.810 3.300 3.150 4.155 ;
        RECT  0.550 3.685 2.810 4.155 ;
        RECT  0.170 3.010 0.550 4.155 ;
        RECT  0.000 3.685 0.170 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.355 0.465 8.220 0.695 ;
        RECT  6.730 3.225 8.220 3.455 ;
        RECT  6.490 2.510 6.730 3.455 ;
        RECT  4.990 3.225 6.490 3.455 ;
        RECT  3.565 2.765 6.060 2.995 ;
        RECT  3.125 0.465 3.355 1.410 ;
        RECT  1.915 1.180 3.125 1.410 ;
        RECT  1.685 0.495 1.915 1.410 ;
        RECT  0.470 1.180 1.685 1.410 ;
        RECT  0.240 0.495 0.470 1.410 ;
    END
END OAI32D2BWP7T

MACRO OAI33D0BWP7T
    CLASS CORE ;
    FOREIGN OAI33D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1340 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 3.045 2.605 3.275 ;
        RECT  1.625 0.930 1.965 1.540 ;
        RECT  0.980 1.310 1.625 1.540 ;
        RECT  0.700 1.310 0.980 3.275 ;
        RECT  0.470 1.310 0.700 1.540 ;
        RECT  0.230 0.860 0.470 1.540 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.770 3.220 2.710 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.770 3.780 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.770 4.900 2.190 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.770 2.165 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.770 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.875 -0.235 5.040 0.235 ;
        RECT  4.495 -0.235 4.875 1.120 ;
        RECT  3.430 -0.235 4.495 0.235 ;
        RECT  3.050 -0.235 3.430 1.080 ;
        RECT  0.000 -0.235 3.050 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.765 3.685 5.040 4.155 ;
        RECT  4.385 3.015 4.765 4.155 ;
        RECT  0.465 3.685 4.385 4.155 ;
        RECT  0.235 3.065 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.855 0.835 4.085 1.540 ;
        RECT  2.645 1.310 3.855 1.540 ;
        RECT  2.415 0.465 2.645 1.540 ;
        RECT  1.245 0.465 2.415 0.695 ;
        RECT  0.905 0.465 1.245 1.080 ;
    END
END OAI33D0BWP7T

MACRO OAI33D1BWP7T
    CLASS CORE ;
    FOREIGN OAI33D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 2.2680 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.980 3.045 2.605 3.275 ;
        RECT  1.625 0.930 1.965 1.345 ;
        RECT  0.980 1.115 1.625 1.345 ;
        RECT  0.700 1.115 0.980 3.275 ;
        RECT  0.470 1.115 0.700 1.345 ;
        RECT  0.230 0.490 0.470 1.345 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.875 1.640 3.220 2.710 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.640 3.780 2.710 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.690 4.900 2.190 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.640 2.165 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.625 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.625 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.815 -0.235 5.040 0.235 ;
        RECT  4.565 -0.235 4.815 1.245 ;
        RECT  3.430 -0.235 4.565 0.235 ;
        RECT  3.050 -0.235 3.430 0.885 ;
        RECT  0.000 -0.235 3.050 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.740 3.685 5.040 4.155 ;
        RECT  4.400 2.535 4.740 4.155 ;
        RECT  0.465 3.685 4.400 4.155 ;
        RECT  0.235 3.065 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.855 0.485 4.085 1.345 ;
        RECT  2.645 1.115 3.855 1.345 ;
        RECT  2.415 0.465 2.645 1.345 ;
        RECT  1.245 0.465 2.415 0.695 ;
        RECT  0.905 0.465 1.245 0.830 ;
    END
END OAI33D1BWP7T

MACRO OAI33D2BWP7T
    CLASS CORE ;
    FOREIGN OAI33D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 3.4024 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.175 0.925 9.405 3.295 ;
        RECT  5.040 0.925 9.175 1.155 ;
        RECT  8.975 3.015 9.175 3.295 ;
        RECT  5.200 2.530 5.430 3.375 ;
        RECT  4.900 2.530 5.200 2.760 ;
        RECT  4.900 0.925 5.040 1.590 ;
        RECT  4.810 0.925 4.900 2.760 ;
        RECT  4.620 1.360 4.810 2.760 ;
        RECT  4.270 2.530 4.620 2.760 ;
        RECT  4.040 2.530 4.270 3.280 ;
        RECT  2.075 3.050 4.040 3.280 ;
        END
    END ZN
    PIN B3
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.820 2.710 2.100 ;
        END
    END B3
    PIN B2
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.910 3.350 2.150 ;
        RECT  2.940 1.360 3.220 2.150 ;
        RECT  1.540 1.360 2.940 1.590 ;
        RECT  1.245 1.360 1.540 2.150 ;
        END
    END B2
    PIN B1
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.810 1.490 4.265 1.725 ;
        RECT  3.580 1.490 3.810 2.710 ;
        RECT  0.980 2.480 3.580 2.710 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.415 1.920 0.700 2.150 ;
        END
    END B1
    PIN A3
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 1.865 8.945 2.205 ;
        RECT  8.540 1.385 8.820 2.710 ;
        RECT  5.510 1.385 8.540 1.615 ;
        RECT  5.280 1.385 5.510 2.025 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.045 1.845 8.275 3.220 ;
        RECT  6.340 2.940 8.045 3.220 ;
        RECT  6.110 1.865 6.340 3.220 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.7848 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.360 2.380 7.750 2.660 ;
        RECT  7.020 1.845 7.360 2.660 ;
        RECT  6.810 2.380 7.020 2.660 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.120 -0.235 9.520 0.235 ;
        RECT  3.780 -0.235 4.120 0.670 ;
        RECT  2.680 -0.235 3.780 0.235 ;
        RECT  2.340 -0.235 2.680 0.670 ;
        RECT  1.240 -0.235 2.340 0.235 ;
        RECT  0.895 -0.235 1.240 0.670 ;
        RECT  0.000 -0.235 0.895 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.350 3.685 9.520 4.155 ;
        RECT  6.990 3.455 7.350 4.155 ;
        RECT  4.730 3.685 6.990 4.155 ;
        RECT  4.500 3.195 4.730 4.155 ;
        RECT  0.465 3.685 4.500 4.155 ;
        RECT  0.235 2.575 0.465 4.155 ;
        RECT  0.000 3.685 0.235 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.580 0.465 9.330 0.695 ;
        RECT  4.350 0.465 4.580 1.130 ;
        RECT  0.465 0.900 4.350 1.130 ;
        RECT  0.235 0.665 0.465 1.130 ;
    END
END OAI33D2BWP7T

MACRO OR2D0BWP7T
    CLASS CORE ;
    FOREIGN OR2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.925 2.660 3.345 ;
        RECT  2.280 0.925 2.380 1.155 ;
        RECT  2.280 3.115 2.380 3.345 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.170 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.535 -0.235 2.800 0.235 ;
        RECT  0.180 -0.235 0.535 0.465 ;
        RECT  0.000 -0.235 0.180 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.865 3.685 2.800 4.155 ;
        RECT  1.520 3.170 1.865 4.155 ;
        RECT  0.000 3.685 1.520 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.025 1.830 2.140 2.170 ;
        RECT  1.785 0.915 2.025 2.940 ;
        RECT  0.940 0.915 1.785 1.145 ;
        RECT  0.510 2.710 1.785 2.940 ;
        RECT  0.270 2.710 0.510 3.420 ;
    END
END OR2D0BWP7T

MACRO OR2D1BWP7T
    CLASS CORE ;
    FOREIGN OR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.465 2.660 3.350 ;
        RECT  2.335 0.465 2.380 1.275 ;
        RECT  2.335 2.380 2.380 3.350 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.735 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 -0.235 2.800 0.235 ;
        RECT  0.140 -0.235 0.550 0.465 ;
        RECT  0.000 -0.235 0.140 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 3.685 2.800 4.155 ;
        RECT  1.505 3.030 1.885 4.155 ;
        RECT  0.000 3.685 1.505 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.020 1.680 2.135 2.020 ;
        RECT  1.780 1.015 2.020 2.800 ;
        RECT  0.940 1.015 1.780 1.245 ;
        RECT  0.505 2.540 1.780 2.800 ;
        RECT  0.275 2.540 0.505 3.350 ;
    END
END OR2D1BWP7T

MACRO OR2D2BWP7T
    CLASS CORE ;
    FOREIGN OR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.665 2.440 2.765 3.250 ;
        RECT  2.380 0.470 2.665 3.250 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.735 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 -0.235 3.920 0.235 ;
        RECT  3.100 -0.235 3.440 1.195 ;
        RECT  2.005 -0.235 3.100 0.235 ;
        RECT  1.655 -0.235 2.005 0.710 ;
        RECT  0.580 -0.235 1.655 0.235 ;
        RECT  0.200 -0.235 0.580 0.710 ;
        RECT  0.000 -0.235 0.200 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.550 3.685 3.920 4.155 ;
        RECT  3.200 2.545 3.550 4.155 ;
        RECT  2.115 3.685 3.200 4.155 ;
        RECT  1.735 2.935 2.115 4.155 ;
        RECT  0.000 3.685 1.735 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.880 0.940 2.140 2.670 ;
        RECT  1.225 0.940 1.880 1.180 ;
        RECT  1.080 2.430 1.880 2.670 ;
        RECT  0.995 0.465 1.225 1.180 ;
        RECT  0.820 2.430 1.080 3.210 ;
        RECT  0.180 2.980 0.820 3.210 ;
    END
END OR2D2BWP7T

MACRO OR2D4BWP7T
    CLASS CORE ;
    FOREIGN OR2D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.535 1.375 5.770 3.220 ;
        RECT  5.505 1.375 5.535 2.780 ;
        RECT  5.275 0.495 5.505 2.780 ;
        RECT  4.870 1.040 5.275 2.780 ;
        RECT  4.065 1.040 4.870 1.390 ;
        RECT  4.325 2.430 4.870 2.780 ;
        RECT  4.095 2.430 4.325 3.240 ;
        RECT  3.835 0.495 4.065 1.390 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 1.660 2.865 2.660 ;
        RECT  0.980 2.380 2.635 2.660 ;
        RECT  0.700 1.660 0.980 2.660 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.660 2.135 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.300 -0.235 6.720 0.235 ;
        RECT  5.920 -0.235 6.300 1.195 ;
        RECT  4.870 -0.235 5.920 0.235 ;
        RECT  4.490 -0.235 4.870 0.785 ;
        RECT  3.440 -0.235 4.490 0.235 ;
        RECT  3.060 -0.235 3.440 0.710 ;
        RECT  2.000 -0.235 3.060 0.235 ;
        RECT  1.620 -0.235 2.000 0.710 ;
        RECT  0.540 -0.235 1.620 0.235 ;
        RECT  0.160 -0.235 0.540 0.710 ;
        RECT  0.000 -0.235 0.160 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 3.685 6.720 4.155 ;
        RECT  6.250 2.245 6.490 4.155 ;
        RECT  5.130 3.685 6.250 4.155 ;
        RECT  4.750 3.060 5.130 4.155 ;
        RECT  3.545 3.685 4.750 4.155 ;
        RECT  3.155 3.350 3.545 4.155 ;
        RECT  0.470 3.685 3.155 4.155 ;
        RECT  0.230 2.245 0.470 4.155 ;
        RECT  0.000 3.685 0.230 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.065 1.040 4.670 1.390 ;
        RECT  4.325 2.430 4.670 2.780 ;
        RECT  4.095 2.430 4.325 3.240 ;
        RECT  3.835 0.495 4.065 1.390 ;
        RECT  3.480 1.755 4.585 1.985 ;
        RECT  3.210 1.040 3.480 3.120 ;
        RECT  2.625 1.040 3.210 1.280 ;
        RECT  1.620 2.890 3.210 3.120 ;
        RECT  2.395 0.465 2.625 1.280 ;
        RECT  1.185 1.040 2.395 1.280 ;
        RECT  0.955 0.465 1.185 1.280 ;
    END
END OR2D4BWP7T

MACRO OR2D8BWP7T
    CLASS CORE ;
    FOREIGN OR2D8BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 5.1192 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 0.495 9.690 3.230 ;
        RECT  8.790 1.040 9.455 2.730 ;
        RECT  8.245 1.040 8.790 1.390 ;
        RECT  8.245 2.380 8.790 2.730 ;
        RECT  8.015 0.495 8.245 1.390 ;
        RECT  8.015 2.380 8.245 3.230 ;
        RECT  6.805 1.040 8.015 1.390 ;
        RECT  6.805 2.380 8.015 2.730 ;
        RECT  6.575 0.495 6.805 1.390 ;
        RECT  6.575 2.380 6.805 3.230 ;
        RECT  5.365 1.040 6.575 1.390 ;
        RECT  5.365 2.380 6.575 2.730 ;
        RECT  5.135 0.495 5.365 1.390 ;
        RECT  5.135 2.380 5.365 3.230 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 1.0098 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.600 4.340 2.710 ;
        RECT  1.540 2.470 4.060 2.710 ;
        RECT  1.200 1.735 1.540 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 1.0098 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.695 3.425 2.150 ;
        RECT  2.380 1.265 2.660 2.150 ;
        RECT  0.685 1.265 2.380 1.505 ;
        RECT  0.455 1.265 0.685 1.940 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.475 -0.235 10.640 0.235 ;
        RECT  10.095 -0.235 10.475 1.250 ;
        RECT  9.045 -0.235 10.095 0.235 ;
        RECT  8.665 -0.235 9.045 0.785 ;
        RECT  7.605 -0.235 8.665 0.235 ;
        RECT  7.225 -0.235 7.605 0.785 ;
        RECT  6.170 -0.235 7.225 0.235 ;
        RECT  5.790 -0.235 6.170 0.785 ;
        RECT  4.730 -0.235 5.790 0.235 ;
        RECT  4.350 -0.235 4.730 0.690 ;
        RECT  3.220 -0.235 4.350 0.235 ;
        RECT  2.880 -0.235 3.220 0.575 ;
        RECT  1.680 -0.235 2.880 0.235 ;
        RECT  1.340 -0.235 1.680 0.925 ;
        RECT  0.000 -0.235 1.340 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.415 3.685 10.640 4.155 ;
        RECT  10.155 2.240 10.415 4.155 ;
        RECT  9.055 3.685 10.155 4.155 ;
        RECT  8.675 2.995 9.055 4.155 ;
        RECT  7.615 3.685 8.675 4.155 ;
        RECT  7.235 2.995 7.615 4.155 ;
        RECT  6.180 3.685 7.235 4.155 ;
        RECT  5.800 2.995 6.180 4.155 ;
        RECT  4.630 3.685 5.800 4.155 ;
        RECT  4.280 3.400 4.630 4.155 ;
        RECT  1.880 3.685 4.280 4.155 ;
        RECT  1.520 3.400 1.880 4.155 ;
        RECT  0.000 3.685 1.520 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.245 1.040 8.590 1.390 ;
        RECT  8.245 2.380 8.590 2.730 ;
        RECT  8.015 0.495 8.245 1.390 ;
        RECT  8.015 2.380 8.245 3.230 ;
        RECT  6.805 1.040 8.015 1.390 ;
        RECT  6.805 2.380 8.015 2.730 ;
        RECT  6.575 0.495 6.805 1.390 ;
        RECT  6.575 2.380 6.805 3.230 ;
        RECT  5.365 1.040 6.575 1.390 ;
        RECT  5.365 2.380 6.575 2.730 ;
        RECT  5.135 0.495 5.365 1.390 ;
        RECT  5.135 2.380 5.365 3.230 ;
        RECT  4.905 1.655 8.470 1.885 ;
        RECT  4.665 1.050 4.905 3.170 ;
        RECT  3.925 1.050 4.665 1.290 ;
        RECT  0.465 2.940 4.665 3.170 ;
        RECT  3.695 0.465 3.925 1.290 ;
        RECT  2.345 0.805 3.695 1.035 ;
        RECT  2.115 0.465 2.345 1.035 ;
        RECT  0.235 2.355 0.465 3.170 ;
    END
END OR2D8BWP7T

MACRO OR2XD1BWP7T
    CLASS CORE ;
    FOREIGN OR2XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 0.495 2.660 3.390 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.590 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.450 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.980 -0.235 3.360 0.235 ;
        RECT  1.600 -0.235 1.980 0.855 ;
        RECT  0.545 -0.235 1.600 0.235 ;
        RECT  0.165 -0.235 0.545 0.930 ;
        RECT  0.000 -0.235 0.165 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 3.685 3.360 4.155 ;
        RECT  1.610 2.940 1.990 4.155 ;
        RECT  0.000 3.685 1.610 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.905 1.110 2.145 2.710 ;
        RECT  1.185 1.110 1.905 1.350 ;
        RECT  0.565 2.470 1.905 2.710 ;
        RECT  0.955 0.495 1.185 1.350 ;
        RECT  0.335 2.470 0.565 3.340 ;
    END
END OR2XD1BWP7T

MACRO OR3D0BWP7T
    CLASS CORE ;
    FOREIGN OR3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.485 3.780 3.345 ;
        RECT  3.190 0.485 3.500 0.725 ;
        RECT  2.900 3.115 3.500 3.345 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.770 0.465 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.190 1.455 1.540 2.150 ;
        RECT  0.700 1.770 1.190 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.770 2.660 2.280 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.805 -0.235 3.920 0.235 ;
        RECT  2.455 -0.235 2.805 0.695 ;
        RECT  1.295 -0.235 2.455 0.235 ;
        RECT  0.930 -0.235 1.295 0.685 ;
        RECT  0.000 -0.235 0.930 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.505 3.685 3.920 4.155 ;
        RECT  2.125 3.235 2.505 4.155 ;
        RECT  0.000 3.685 2.125 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.910 0.955 3.140 2.885 ;
        RECT  1.985 0.955 2.910 1.215 ;
        RECT  1.670 2.645 2.910 2.885 ;
        RECT  1.755 0.480 1.985 1.215 ;
        RECT  0.465 0.955 1.755 1.215 ;
        RECT  1.440 2.645 1.670 3.285 ;
        RECT  0.180 3.055 1.440 3.285 ;
        RECT  0.235 0.480 0.465 1.215 ;
    END
END OR3D0BWP7T

MACRO OR3D1BWP7T
    CLASS CORE ;
    FOREIGN OR3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2192 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.495 3.780 3.080 ;
        RECT  3.280 0.495 3.500 1.305 ;
        RECT  2.905 2.850 3.500 3.080 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.730 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.150 ;
        RECT  1.180 1.210 1.260 1.480 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.145 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.800 -0.235 3.920 0.235 ;
        RECT  2.455 -0.235 2.800 0.505 ;
        RECT  1.280 -0.235 2.455 0.235 ;
        RECT  0.935 -0.235 1.280 0.505 ;
        RECT  0.000 -0.235 0.935 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 3.685 3.920 4.155 ;
        RECT  2.130 2.850 2.510 4.155 ;
        RECT  0.000 3.685 2.130 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.800 0.735 3.050 2.620 ;
        RECT  1.985 0.735 2.800 0.965 ;
        RECT  0.475 2.380 2.800 2.620 ;
        RECT  1.755 0.465 1.985 0.965 ;
        RECT  0.465 0.735 1.755 0.965 ;
        RECT  0.225 2.380 0.475 3.335 ;
        RECT  0.235 0.465 0.465 0.965 ;
    END
END OR3D1BWP7T

MACRO OR3D2BWP7T
    CLASS CORE ;
    FOREIGN OR3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 1.065 3.780 2.150 ;
        RECT  3.500 0.495 3.525 2.150 ;
        RECT  3.295 0.495 3.500 1.305 ;
        RECT  3.410 1.890 3.500 2.150 ;
        RECT  3.170 1.890 3.410 3.145 ;
        RECT  2.880 2.915 3.170 3.145 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.680 0.980 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 1.210 1.550 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.210 2.125 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.250 -0.235 4.480 0.235 ;
        RECT  4.015 -0.235 4.250 1.250 ;
        RECT  2.840 -0.235 4.015 0.235 ;
        RECT  2.470 -0.235 2.840 0.490 ;
        RECT  1.300 -0.235 2.470 0.235 ;
        RECT  0.955 -0.235 1.300 0.490 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.885 3.685 4.480 4.155 ;
        RECT  3.655 2.535 3.885 4.155 ;
        RECT  2.460 3.685 3.655 4.155 ;
        RECT  2.100 2.925 2.460 4.155 ;
        RECT  0.000 3.685 2.100 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.710 0.720 2.940 2.620 ;
        RECT  2.005 0.720 2.710 0.980 ;
        RECT  0.490 2.380 2.710 2.620 ;
        RECT  1.775 0.480 2.005 0.980 ;
        RECT  0.485 0.720 1.775 0.980 ;
        RECT  0.250 2.380 0.490 3.245 ;
        RECT  0.255 0.480 0.485 0.980 ;
    END
END OR3D2BWP7T

MACRO OR3D4BWP7T
    CLASS CORE ;
    FOREIGN OR3D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.095 0.475 6.330 3.245 ;
        RECT  5.430 1.080 6.095 2.690 ;
        RECT  4.885 1.080 5.430 1.430 ;
        RECT  4.885 2.420 5.430 2.690 ;
        RECT  4.655 0.475 4.885 1.430 ;
        RECT  4.655 2.420 4.885 3.245 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.370 1.780 2.710 2.100 ;
        RECT  1.770 1.820 2.370 2.100 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.070 1.155 3.410 1.540 ;
        RECT  1.530 1.260 3.070 1.540 ;
        RECT  1.300 1.260 1.530 2.065 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 1.725 3.925 2.495 ;
        RECT  3.195 2.255 3.695 2.495 ;
        RECT  2.955 2.255 3.195 2.710 ;
        RECT  0.450 2.480 2.955 2.710 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.100 -0.235 7.280 0.235 ;
        RECT  6.760 -0.235 7.100 1.195 ;
        RECT  5.660 -0.235 6.760 0.235 ;
        RECT  5.320 -0.235 5.660 0.850 ;
        RECT  4.180 -0.235 5.320 0.235 ;
        RECT  3.840 -0.235 4.180 0.465 ;
        RECT  2.105 -0.235 3.840 0.235 ;
        RECT  1.765 -0.235 2.105 0.465 ;
        RECT  0.575 -0.235 1.765 0.235 ;
        RECT  0.235 -0.235 0.575 1.190 ;
        RECT  0.000 -0.235 0.235 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.100 3.685 7.280 4.155 ;
        RECT  6.760 2.565 7.100 4.155 ;
        RECT  5.660 3.685 6.760 4.155 ;
        RECT  5.320 2.920 5.660 4.155 ;
        RECT  4.165 3.685 5.320 4.155 ;
        RECT  3.935 3.195 4.165 4.155 ;
        RECT  0.615 3.685 3.935 4.155 ;
        RECT  0.275 3.130 0.615 4.155 ;
        RECT  0.000 3.685 0.275 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.885 1.080 5.230 1.430 ;
        RECT  4.885 2.420 5.230 2.690 ;
        RECT  4.655 0.475 4.885 1.430 ;
        RECT  4.655 2.420 4.885 3.245 ;
        RECT  4.425 1.715 5.170 1.945 ;
        RECT  4.185 0.695 4.425 2.965 ;
        RECT  1.005 0.695 4.185 0.925 ;
        RECT  3.665 2.725 4.185 2.965 ;
        RECT  3.425 2.725 3.665 3.270 ;
        RECT  2.255 3.040 3.425 3.270 ;
    END
END OR3D4BWP7T

MACRO OR3XD1BWP7T
    CLASS CORE ;
    FOREIGN OR3XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 0.580 3.780 2.820 ;
        RECT  3.125 0.580 3.500 0.810 ;
        RECT  3.410 2.580 3.500 2.820 ;
        RECT  3.180 2.580 3.410 3.390 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.660 0.450 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.660 1.540 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.660 2.665 2.710 ;
        RECT  2.230 1.660 2.380 2.000 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 -0.235 3.920 0.235 ;
        RECT  2.390 -0.235 2.770 0.810 ;
        RECT  1.330 -0.235 2.390 0.235 ;
        RECT  0.950 -0.235 1.330 0.810 ;
        RECT  0.000 -0.235 0.950 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.680 3.685 3.920 4.155 ;
        RECT  2.300 3.025 2.680 4.155 ;
        RECT  0.000 3.685 2.300 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.940 1.040 3.170 2.000 ;
        RECT  2.000 1.040 2.940 1.290 ;
        RECT  1.970 1.040 2.000 3.170 ;
        RECT  1.770 0.480 1.970 3.170 ;
        RECT  1.740 0.480 1.770 1.290 ;
        RECT  0.300 2.940 1.770 3.170 ;
        RECT  0.530 1.040 1.740 1.290 ;
        RECT  0.300 0.480 0.530 1.290 ;
    END
END OR3XD1BWP7T

MACRO OR4D0BWP7T
    CLASS CORE ;
    FOREIGN OR4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.625 4.340 3.345 ;
        RECT  3.925 0.625 4.060 0.855 ;
        RECT  3.940 3.115 4.060 3.345 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        RECT  0.580 1.630 0.700 1.970 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.595 2.200 1.825 ;
        RECT  1.820 1.595 2.100 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.770 3.220 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.520 -0.235 4.480 0.235 ;
        RECT  3.180 -0.235 3.520 0.490 ;
        RECT  2.015 -0.235 3.180 0.235 ;
        RECT  1.630 -0.235 2.015 0.490 ;
        RECT  0.555 -0.235 1.630 0.235 ;
        RECT  0.175 -0.235 0.555 0.825 ;
        RECT  0.000 -0.235 0.175 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.355 3.685 4.480 4.155 ;
        RECT  2.970 3.450 3.355 4.155 ;
        RECT  0.000 3.685 2.970 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.460 0.720 3.690 3.220 ;
        RECT  2.705 0.720 3.460 0.960 ;
        RECT  0.280 2.990 3.460 3.220 ;
        RECT  2.475 0.540 2.705 0.960 ;
        RECT  1.185 0.720 2.475 0.960 ;
        RECT  0.955 0.540 1.185 0.960 ;
    END
END OR4D0BWP7T

MACRO OR4D1BWP7T
    CLASS CORE ;
    FOREIGN OR4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.495 4.340 3.070 ;
        RECT  3.980 0.495 4.060 1.305 ;
        RECT  3.555 2.840 4.060 3.070 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.685 0.980 2.710 ;
        RECT  0.580 1.685 0.700 2.025 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.440 1.540 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.385 2.150 1.725 ;
        RECT  1.820 1.385 2.100 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.510 -0.235 4.480 0.235 ;
        RECT  3.160 -0.235 3.510 0.685 ;
        RECT  2.060 -0.235 3.160 0.235 ;
        RECT  1.660 -0.235 2.060 0.685 ;
        RECT  0.610 -0.235 1.660 0.235 ;
        RECT  0.230 -0.235 0.610 0.750 ;
        RECT  0.000 -0.235 0.230 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.170 3.685 4.480 4.155 ;
        RECT  2.790 2.840 3.170 4.155 ;
        RECT  0.000 3.685 2.790 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.455 0.915 3.685 2.610 ;
        RECT  2.745 0.915 3.455 1.155 ;
        RECT  2.560 2.380 3.455 2.610 ;
        RECT  2.395 0.515 2.745 1.155 ;
        RECT  2.330 2.380 2.560 3.170 ;
        RECT  1.295 0.915 2.395 1.155 ;
        RECT  0.280 2.940 2.330 3.170 ;
        RECT  0.950 0.520 1.295 1.155 ;
    END
END OR4D1BWP7T

MACRO OR4D2BWP7T
    CLASS CORE ;
    FOREIGN OR4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 1.210 4.340 2.720 ;
        RECT  4.060 1.210 4.085 3.290 ;
        RECT  4.005 1.210 4.060 1.450 ;
        RECT  3.855 2.390 4.060 3.290 ;
        RECT  3.775 0.495 4.005 1.450 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.140 1.210 0.465 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.240 1.680 1.540 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.680 2.140 3.270 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.3366 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 1.770 2.925 2.010 ;
        RECT  2.380 1.770 2.660 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.790 -0.235 5.040 0.235 ;
        RECT  4.435 -0.235 4.790 0.730 ;
        RECT  3.315 -0.235 4.435 0.235 ;
        RECT  2.940 -0.235 3.315 0.480 ;
        RECT  0.525 -0.235 2.940 0.235 ;
        RECT  0.140 -0.235 0.525 0.825 ;
        RECT  0.000 -0.235 0.140 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.810 3.685 5.040 4.155 ;
        RECT  4.575 2.240 4.810 4.155 ;
        RECT  3.280 3.685 4.575 4.155 ;
        RECT  2.940 2.585 3.280 4.155 ;
        RECT  0.000 3.685 2.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.390 1.775 3.830 2.005 ;
        RECT  3.160 1.120 3.390 2.005 ;
        RECT  2.505 1.120 3.160 1.400 ;
        RECT  2.275 0.595 2.505 1.400 ;
        RECT  1.010 0.595 2.275 0.825 ;
        RECT  0.770 0.595 1.010 2.730 ;
        RECT  0.555 2.450 0.770 2.730 ;
        RECT  0.325 2.450 0.555 3.320 ;
    END
END OR4D2BWP7T

MACRO OR4D4BWP7T
    CLASS CORE ;
    FOREIGN OR4D4BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.960 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 2.5596 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.775 0.465 8.010 3.260 ;
        RECT  7.110 1.070 7.775 2.570 ;
        RECT  6.565 1.070 7.110 1.420 ;
        RECT  6.565 2.220 7.110 2.570 ;
        RECT  6.335 0.465 6.565 1.420 ;
        RECT  6.335 2.220 6.565 3.300 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.670 1.260 4.390 1.540 ;
        RECT  3.440 1.260 3.670 2.010 ;
        RECT  3.125 1.780 3.440 2.010 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.130 1.780 4.240 2.010 ;
        RECT  3.900 1.780 4.130 2.535 ;
        RECT  2.660 2.305 3.900 2.535 ;
        RECT  2.430 1.770 2.660 2.535 ;
        RECT  1.820 1.770 2.430 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.730 1.780 4.910 2.010 ;
        RECT  4.500 1.780 4.730 2.995 ;
        RECT  1.540 2.765 4.500 2.995 ;
        RECT  1.250 1.670 1.540 2.995 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.6732 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.295 0.700 5.525 2.000 ;
        RECT  3.210 0.700 5.295 0.930 ;
        RECT  2.980 0.700 3.210 1.440 ;
        RECT  0.980 1.210 2.980 1.440 ;
        RECT  0.700 1.210 0.980 2.190 ;
        RECT  0.580 1.660 0.700 2.000 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.815 -0.235 8.960 0.235 ;
        RECT  8.435 -0.235 8.815 1.200 ;
        RECT  7.375 -0.235 8.435 0.235 ;
        RECT  6.995 -0.235 7.375 0.825 ;
        RECT  5.860 -0.235 6.995 0.235 ;
        RECT  5.520 -0.235 5.860 0.465 ;
        RECT  3.565 -0.235 5.520 0.235 ;
        RECT  3.225 -0.235 3.565 0.465 ;
        RECT  2.045 -0.235 3.225 0.235 ;
        RECT  1.705 -0.235 2.045 0.465 ;
        RECT  0.525 -0.235 1.705 0.235 ;
        RECT  0.185 -0.235 0.525 0.465 ;
        RECT  0.000 -0.235 0.185 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.810 3.685 8.960 4.155 ;
        RECT  8.430 2.565 8.810 4.155 ;
        RECT  7.355 3.685 8.430 4.155 ;
        RECT  6.975 2.880 7.355 4.155 ;
        RECT  5.860 3.685 6.975 4.155 ;
        RECT  5.520 3.455 5.860 4.155 ;
        RECT  0.540 3.685 5.520 4.155 ;
        RECT  0.310 3.195 0.540 4.155 ;
        RECT  0.000 3.685 0.310 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.565 1.070 6.910 1.420 ;
        RECT  6.565 2.220 6.910 2.570 ;
        RECT  6.335 0.465 6.565 1.420 ;
        RECT  6.335 2.220 6.565 3.300 ;
        RECT  6.105 1.715 6.880 1.945 ;
        RECT  5.875 1.020 6.105 3.130 ;
        RECT  5.240 2.890 5.875 3.130 ;
        RECT  5.000 2.890 5.240 3.455 ;
        RECT  1.020 3.225 5.000 3.455 ;
        RECT  0.350 0.695 2.520 0.925 ;
        RECT  0.790 2.445 1.020 3.455 ;
        RECT  0.350 2.445 0.790 2.675 ;
        RECT  0.120 0.695 0.350 2.675 ;
        RECT  2.520 0.575 2.750 0.925 ;
    END
END OR4D4BWP7T

MACRO OR4XD1BWP7T
    CLASS CORE ;
    FOREIGN OR4XD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 0.640 4.340 3.175 ;
        RECT  3.835 0.640 4.060 0.870 ;
        RECT  3.595 2.945 4.060 3.175 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.420 1.715 0.845 1.945 ;
        RECT  0.140 1.715 0.420 2.710 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.660 1.540 2.710 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.660 2.150 2.000 ;
        RECT  1.820 1.660 2.100 2.710 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.770 3.220 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 -0.235 4.480 0.235 ;
        RECT  3.115 -0.235 3.455 0.810 ;
        RECT  2.015 -0.235 3.115 0.235 ;
        RECT  1.675 -0.235 2.015 0.810 ;
        RECT  0.560 -0.235 1.675 0.235 ;
        RECT  0.220 -0.235 0.560 1.200 ;
        RECT  0.000 -0.235 0.220 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.240 3.685 4.480 4.155 ;
        RECT  2.860 2.900 3.240 4.155 ;
        RECT  0.000 3.685 2.860 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.450 1.040 3.680 2.670 ;
        RECT  2.680 1.040 3.450 1.320 ;
        RECT  2.605 2.430 3.450 2.670 ;
        RECT  2.450 0.485 2.680 1.320 ;
        RECT  2.365 2.430 2.605 3.295 ;
        RECT  1.225 1.040 2.450 1.320 ;
        RECT  0.265 3.065 2.365 3.295 ;
        RECT  0.995 0.490 1.225 1.320 ;
    END
END OR4XD1BWP7T

MACRO SDFCND0BWP7T
    CLASS CORE ;
    FOREIGN SDFCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.150 15.540 2.560 ;
        RECT  15.125 1.150 15.260 1.380 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.585 15.125 1.380 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.590 16.660 2.705 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.600 3.780 2.710 ;
        RECT  3.380 1.600 3.500 1.940 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.470 1.615 4.620 1.955 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.225 11.925 3.455 ;
        RECT  10.805 2.730 11.035 3.455 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.885 ;
        RECT  12.255 -0.235 15.560 0.235 ;
        RECT  11.915 -0.235 12.255 0.465 ;
        RECT  8.955 -0.235 11.915 0.235 ;
        RECT  8.615 -0.235 8.955 1.100 ;
        RECT  4.145 -0.235 8.615 0.235 ;
        RECT  3.805 -0.235 4.145 0.465 ;
        RECT  1.240 -0.235 3.805 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.820 3.685 16.800 4.155 ;
        RECT  15.480 3.455 15.820 4.155 ;
        RECT  14.640 3.685 15.480 4.155 ;
        RECT  14.300 3.455 14.640 4.155 ;
        RECT  13.110 3.685 14.300 4.155 ;
        RECT  12.770 3.190 13.110 4.155 ;
        RECT  10.575 3.685 12.770 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.975 3.685 10.235 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  14.575 2.790 15.855 3.020 ;
        RECT  12.850 0.465 14.660 0.695 ;
        RECT  14.345 0.990 14.575 3.020 ;
        RECT  13.455 0.990 14.345 1.220 ;
        RECT  13.820 2.555 14.345 2.785 ;
        RECT  13.835 1.565 14.065 2.325 ;
        RECT  13.015 2.095 13.835 2.325 ;
        RECT  13.590 2.555 13.820 3.420 ;
        RECT  13.225 0.990 13.455 1.865 ;
        RECT  12.280 1.635 13.225 1.865 ;
        RECT  12.785 2.095 13.015 2.960 ;
        RECT  12.620 0.465 12.850 1.220 ;
        RECT  11.495 2.730 12.785 2.960 ;
        RECT  12.000 0.990 12.620 1.220 ;
        RECT  12.000 2.270 12.270 2.500 ;
        RECT  11.770 0.990 12.000 2.500 ;
        RECT  11.015 0.990 11.770 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.755 1.330 9.810 1.560 ;
        RECT  9.525 0.870 9.755 1.560 ;
        RECT  8.805 1.330 9.525 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.280 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  7.100 0.935 7.280 2.230 ;
        RECT  7.050 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.050 3.085 ;
        RECT  6.380 0.780 6.560 2.505 ;
        RECT  6.330 0.780 6.380 3.225 ;
        RECT  6.150 2.275 6.330 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.850 1.615 6.095 1.955 ;
        RECT  5.620 0.760 5.850 2.765 ;
        RECT  5.390 2.535 5.620 2.765 ;
        RECT  5.160 0.975 5.390 1.970 ;
        RECT  4.240 0.975 5.160 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.440 ;
        RECT  2.600 3.210 3.315 3.440 ;
        RECT  3.095 0.475 3.200 1.285 ;
        RECT  2.970 0.475 3.095 2.925 ;
        RECT  2.865 1.090 2.970 2.925 ;
        RECT  2.480 1.075 2.600 3.440 ;
        RECT  2.370 0.465 2.480 3.440 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFCND0BWP7T

MACRO SDFCND1BWP7T
    CLASS CORE ;
    FOREIGN SDFCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.9672 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.075 15.540 2.560 ;
        RECT  15.125 1.075 15.260 1.305 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.480 15.125 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.470 16.660 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.600 3.780 2.710 ;
        RECT  3.380 1.600 3.500 1.940 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.470 1.615 4.620 1.955 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.225 11.925 3.455 ;
        RECT  10.805 2.730 11.035 3.455 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.810 ;
        RECT  12.255 -0.235 15.560 0.235 ;
        RECT  11.915 -0.235 12.255 0.465 ;
        RECT  8.955 -0.235 11.915 0.235 ;
        RECT  8.615 -0.235 8.955 1.100 ;
        RECT  4.145 -0.235 8.615 0.235 ;
        RECT  3.805 -0.235 4.145 0.465 ;
        RECT  1.240 -0.235 3.805 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 3.685 16.800 4.155 ;
        RECT  15.560 3.250 15.900 4.155 ;
        RECT  14.640 3.685 15.560 4.155 ;
        RECT  14.300 3.455 14.640 4.155 ;
        RECT  13.110 3.685 14.300 4.155 ;
        RECT  12.770 3.190 13.110 4.155 ;
        RECT  10.575 3.685 12.770 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.975 3.685 10.235 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  14.575 2.790 15.855 3.020 ;
        RECT  12.850 0.465 14.660 0.695 ;
        RECT  14.345 1.020 14.575 3.020 ;
        RECT  13.455 1.020 14.345 1.250 ;
        RECT  13.820 2.565 14.345 2.795 ;
        RECT  13.835 1.565 14.065 2.260 ;
        RECT  13.015 2.030 13.835 2.260 ;
        RECT  13.590 2.565 13.820 3.375 ;
        RECT  13.225 1.020 13.455 1.760 ;
        RECT  12.280 1.530 13.225 1.760 ;
        RECT  12.785 2.030 13.015 2.960 ;
        RECT  12.620 0.465 12.850 1.220 ;
        RECT  11.495 2.730 12.785 2.960 ;
        RECT  12.000 0.990 12.620 1.220 ;
        RECT  12.000 2.270 12.270 2.500 ;
        RECT  11.770 0.990 12.000 2.500 ;
        RECT  11.015 0.990 11.770 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.755 1.330 9.810 1.560 ;
        RECT  9.525 0.870 9.755 1.560 ;
        RECT  8.805 1.330 9.525 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.280 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  7.100 0.935 7.280 2.230 ;
        RECT  7.050 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.050 3.085 ;
        RECT  6.380 0.745 6.560 2.505 ;
        RECT  6.330 0.745 6.380 3.225 ;
        RECT  6.150 2.275 6.330 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.850 1.615 6.095 1.955 ;
        RECT  5.620 0.720 5.850 2.765 ;
        RECT  5.390 2.535 5.620 2.765 ;
        RECT  5.160 0.975 5.390 1.970 ;
        RECT  4.240 0.975 5.160 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.440 ;
        RECT  2.600 3.210 3.315 3.440 ;
        RECT  3.095 0.475 3.200 1.285 ;
        RECT  2.970 0.475 3.095 2.925 ;
        RECT  2.865 1.090 2.970 2.925 ;
        RECT  2.480 1.075 2.600 3.440 ;
        RECT  2.370 0.465 2.480 3.440 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFCND1BWP7T

MACRO SDFCND2BWP7T
    CLASS CORE ;
    FOREIGN SDFCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.240 0.465 15.585 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 1.055 17.220 2.690 ;
        RECT  16.940 0.465 16.965 3.310 ;
        RECT  16.730 0.465 16.940 1.285 ;
        RECT  16.735 2.460 16.940 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.600 3.780 2.710 ;
        RECT  3.380 1.600 3.500 1.940 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.470 1.615 4.620 1.955 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.190 11.765 3.420 ;
        RECT  10.805 2.730 11.035 3.420 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 -0.235 17.920 0.235 ;
        RECT  17.455 -0.235 17.685 1.245 ;
        RECT  16.300 -0.235 17.455 0.235 ;
        RECT  15.960 -0.235 16.300 1.180 ;
        RECT  14.820 -0.235 15.960 0.235 ;
        RECT  14.480 -0.235 14.820 0.465 ;
        RECT  12.890 -0.235 14.480 0.235 ;
        RECT  12.550 -0.235 12.890 0.465 ;
        RECT  8.955 -0.235 12.550 0.235 ;
        RECT  8.615 -0.235 8.955 1.100 ;
        RECT  4.145 -0.235 8.615 0.235 ;
        RECT  3.805 -0.235 4.145 0.465 ;
        RECT  1.240 -0.235 3.805 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 3.685 17.920 4.155 ;
        RECT  17.455 2.255 17.685 4.155 ;
        RECT  16.300 3.685 17.455 4.155 ;
        RECT  15.960 3.250 16.300 4.155 ;
        RECT  14.705 3.685 15.960 4.155 ;
        RECT  14.365 3.250 14.705 4.155 ;
        RECT  13.105 3.685 14.365 4.155 ;
        RECT  12.765 3.190 13.105 4.155 ;
        RECT  10.575 3.685 12.765 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.975 3.685 10.235 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.255 1.600 16.485 3.020 ;
        RECT  14.480 2.790 16.255 3.020 ;
        RECT  14.770 0.695 15.000 1.940 ;
        RECT  12.075 0.695 14.770 0.925 ;
        RECT  14.250 1.155 14.480 3.020 ;
        RECT  13.035 1.155 14.250 1.385 ;
        RECT  13.825 2.540 14.250 2.770 ;
        RECT  13.720 1.670 13.950 2.260 ;
        RECT  13.595 2.540 13.825 3.370 ;
        RECT  13.055 2.030 13.720 2.260 ;
        RECT  12.825 2.030 13.055 2.960 ;
        RECT  12.805 1.155 13.035 1.750 ;
        RECT  11.495 2.730 12.825 2.960 ;
        RECT  12.305 1.520 12.805 1.750 ;
        RECT  12.075 2.270 12.270 2.500 ;
        RECT  11.845 0.465 12.075 2.500 ;
        RECT  10.970 0.990 11.845 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.655 1.615 11.265 1.845 ;
        RECT  10.425 0.985 10.655 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.425 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.755 1.330 9.810 1.560 ;
        RECT  9.525 0.870 9.755 1.560 ;
        RECT  8.805 1.330 9.525 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.280 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  7.100 0.935 7.280 2.230 ;
        RECT  7.050 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.050 3.085 ;
        RECT  6.380 0.795 6.560 2.505 ;
        RECT  6.330 0.795 6.380 3.225 ;
        RECT  6.150 2.275 6.330 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.850 1.615 6.095 1.955 ;
        RECT  5.620 0.735 5.850 2.765 ;
        RECT  5.390 2.535 5.620 2.765 ;
        RECT  5.160 0.975 5.390 1.970 ;
        RECT  4.240 0.975 5.160 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.440 ;
        RECT  2.600 3.210 3.315 3.440 ;
        RECT  3.095 0.475 3.200 1.285 ;
        RECT  2.970 0.475 3.095 2.925 ;
        RECT  2.865 1.090 2.970 2.925 ;
        RECT  2.480 1.075 2.600 3.440 ;
        RECT  2.370 0.465 2.480 3.440 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFCND2BWP7T

MACRO SDFCNQD0BWP7T
    CLASS CORE ;
    FOREIGN SDFCNQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.210 0.655 15.540 3.400 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.600 3.780 2.710 ;
        RECT  3.380 1.600 3.500 1.940 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.470 1.615 4.620 1.955 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.225 11.925 3.455 ;
        RECT  10.805 2.730 11.035 3.455 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.725 -0.235 15.680 0.235 ;
        RECT  14.495 -0.235 14.725 1.005 ;
        RECT  12.285 -0.235 14.495 0.235 ;
        RECT  11.945 -0.235 12.285 0.465 ;
        RECT  8.955 -0.235 11.945 0.235 ;
        RECT  8.615 -0.235 8.955 1.100 ;
        RECT  4.145 -0.235 8.615 0.235 ;
        RECT  3.805 -0.235 4.145 0.465 ;
        RECT  1.240 -0.235 3.805 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.745 3.685 15.680 4.155 ;
        RECT  14.405 3.115 14.745 4.155 ;
        RECT  13.110 3.685 14.405 4.155 ;
        RECT  12.770 3.190 13.110 4.155 ;
        RECT  10.575 3.685 12.770 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.975 3.685 10.235 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.235 1.600 14.965 1.940 ;
        RECT  14.005 0.990 14.235 2.795 ;
        RECT  13.980 0.990 14.005 1.220 ;
        RECT  13.880 2.565 14.005 2.795 ;
        RECT  13.750 0.465 13.980 1.220 ;
        RECT  13.650 2.565 13.880 3.375 ;
        RECT  13.060 0.990 13.750 1.220 ;
        RECT  13.510 1.565 13.740 2.260 ;
        RECT  13.015 2.030 13.510 2.260 ;
        RECT  12.830 0.990 13.060 1.760 ;
        RECT  12.785 2.030 13.015 2.960 ;
        RECT  12.280 1.530 12.830 1.760 ;
        RECT  11.495 2.730 12.785 2.960 ;
        RECT  12.005 0.990 12.270 1.220 ;
        RECT  12.005 2.270 12.270 2.500 ;
        RECT  11.775 0.990 12.005 2.500 ;
        RECT  11.015 0.990 11.775 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.755 1.330 9.810 1.560 ;
        RECT  9.525 0.870 9.755 1.560 ;
        RECT  8.805 1.330 9.525 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.280 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  7.100 0.935 7.280 2.230 ;
        RECT  7.050 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.050 3.085 ;
        RECT  6.380 0.465 6.560 2.505 ;
        RECT  6.330 0.465 6.380 3.225 ;
        RECT  6.150 2.275 6.330 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.850 1.615 6.095 1.955 ;
        RECT  5.620 0.920 5.850 2.765 ;
        RECT  5.390 2.535 5.620 2.765 ;
        RECT  5.160 0.975 5.390 1.970 ;
        RECT  4.240 0.975 5.160 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.440 ;
        RECT  2.600 3.210 3.315 3.440 ;
        RECT  3.095 0.475 3.200 1.285 ;
        RECT  2.970 0.475 3.095 2.925 ;
        RECT  2.865 1.090 2.970 2.925 ;
        RECT  2.480 1.075 2.600 3.440 ;
        RECT  2.370 0.465 2.480 3.440 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFCNQD0BWP7T

MACRO SDFCNQD1BWP7T
    CLASS CORE ;
    FOREIGN SDFCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.210 0.470 15.540 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.600 3.780 2.710 ;
        RECT  3.380 1.600 3.500 1.940 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.470 1.615 4.620 1.955 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.225 11.925 3.455 ;
        RECT  10.805 2.730 11.035 3.455 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.725 -0.235 15.680 0.235 ;
        RECT  14.495 -0.235 14.725 1.290 ;
        RECT  12.285 -0.235 14.495 0.235 ;
        RECT  11.945 -0.235 12.285 0.465 ;
        RECT  8.955 -0.235 11.945 0.235 ;
        RECT  8.615 -0.235 8.955 1.100 ;
        RECT  4.145 -0.235 8.615 0.235 ;
        RECT  3.805 -0.235 4.145 0.465 ;
        RECT  1.240 -0.235 3.805 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.690 3.685 15.680 4.155 ;
        RECT  14.460 2.255 14.690 4.155 ;
        RECT  13.110 3.685 14.460 4.155 ;
        RECT  12.770 3.190 13.110 4.155 ;
        RECT  10.575 3.685 12.770 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.975 3.685 10.235 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.200 1.600 14.965 1.940 ;
        RECT  13.980 0.990 14.200 2.795 ;
        RECT  13.970 0.465 13.980 2.795 ;
        RECT  13.750 0.465 13.970 1.220 ;
        RECT  13.880 2.565 13.970 2.795 ;
        RECT  13.650 2.565 13.880 3.375 ;
        RECT  13.060 0.990 13.750 1.220 ;
        RECT  13.510 1.565 13.740 2.260 ;
        RECT  13.015 2.030 13.510 2.260 ;
        RECT  12.830 0.990 13.060 1.760 ;
        RECT  12.785 2.030 13.015 2.960 ;
        RECT  12.280 1.530 12.830 1.760 ;
        RECT  11.495 2.730 12.785 2.960 ;
        RECT  12.005 0.990 12.270 1.220 ;
        RECT  12.005 2.270 12.270 2.500 ;
        RECT  11.775 0.990 12.005 2.500 ;
        RECT  11.015 0.990 11.775 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.755 1.330 9.810 1.560 ;
        RECT  9.525 0.870 9.755 1.560 ;
        RECT  8.805 1.330 9.525 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.280 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  7.100 0.935 7.280 2.230 ;
        RECT  7.050 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.050 3.085 ;
        RECT  6.380 0.465 6.560 2.505 ;
        RECT  6.330 0.465 6.380 3.225 ;
        RECT  6.150 2.275 6.330 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.850 1.615 6.095 1.955 ;
        RECT  5.620 0.920 5.850 2.765 ;
        RECT  5.390 2.535 5.620 2.765 ;
        RECT  5.160 0.975 5.390 1.970 ;
        RECT  4.240 0.975 5.160 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.440 ;
        RECT  2.600 3.210 3.315 3.440 ;
        RECT  3.095 0.475 3.200 1.285 ;
        RECT  2.970 0.475 3.095 2.925 ;
        RECT  2.865 1.090 2.970 2.925 ;
        RECT  2.480 1.075 2.600 3.440 ;
        RECT  2.370 0.465 2.480 3.440 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFCNQD1BWP7T

MACRO SDFCNQD2BWP7T
    CLASS CORE ;
    FOREIGN SDFCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.065 15.540 2.730 ;
        RECT  15.260 0.470 15.285 3.310 ;
        RECT  15.050 0.470 15.260 1.295 ;
        RECT  15.055 2.500 15.260 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.600 3.780 2.710 ;
        RECT  3.380 1.600 3.500 1.940 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.470 1.615 4.620 1.955 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.225 11.765 3.455 ;
        RECT  10.805 2.730 11.035 3.455 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.235 ;
        RECT  14.620 -0.235 15.775 0.235 ;
        RECT  14.280 -0.235 14.620 0.755 ;
        RECT  12.185 -0.235 14.280 0.235 ;
        RECT  11.845 -0.235 12.185 0.465 ;
        RECT  8.955 -0.235 11.845 0.235 ;
        RECT  8.615 -0.235 8.955 1.100 ;
        RECT  4.145 -0.235 8.615 0.235 ;
        RECT  3.805 -0.235 4.145 0.465 ;
        RECT  1.240 -0.235 3.805 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.255 16.005 4.155 ;
        RECT  14.615 3.685 15.775 4.155 ;
        RECT  14.275 3.090 14.615 4.155 ;
        RECT  13.110 3.685 14.275 4.155 ;
        RECT  12.770 3.190 13.110 4.155 ;
        RECT  10.575 3.685 12.770 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.975 3.685 10.235 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.550 1.600 14.950 1.940 ;
        RECT  14.320 0.990 14.550 2.795 ;
        RECT  13.865 0.990 14.320 1.220 ;
        RECT  13.835 2.565 14.320 2.795 ;
        RECT  13.635 0.465 13.865 1.220 ;
        RECT  13.635 1.565 13.865 2.260 ;
        RECT  13.605 2.565 13.835 3.375 ;
        RECT  13.005 0.990 13.635 1.220 ;
        RECT  13.015 2.030 13.635 2.260 ;
        RECT  12.785 2.030 13.015 2.960 ;
        RECT  12.775 0.990 13.005 1.760 ;
        RECT  11.495 2.730 12.785 2.960 ;
        RECT  12.230 1.530 12.775 1.760 ;
        RECT  11.985 2.270 12.270 2.500 ;
        RECT  11.985 0.990 12.170 1.220 ;
        RECT  11.755 0.990 11.985 2.500 ;
        RECT  11.015 0.990 11.755 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.755 1.330 9.810 1.560 ;
        RECT  9.525 0.870 9.755 1.560 ;
        RECT  8.805 1.330 9.525 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.280 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  7.100 0.935 7.280 2.230 ;
        RECT  7.050 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.050 3.085 ;
        RECT  6.380 0.465 6.560 2.505 ;
        RECT  6.330 0.465 6.380 3.225 ;
        RECT  6.150 2.275 6.330 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.850 1.615 6.095 1.955 ;
        RECT  5.620 0.920 5.850 2.765 ;
        RECT  5.390 2.535 5.620 2.765 ;
        RECT  5.160 0.975 5.390 1.970 ;
        RECT  4.240 0.975 5.160 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.440 ;
        RECT  2.600 3.210 3.315 3.440 ;
        RECT  3.095 0.475 3.200 1.285 ;
        RECT  2.970 0.475 3.095 2.925 ;
        RECT  2.865 1.090 2.970 2.925 ;
        RECT  2.480 1.075 2.600 3.440 ;
        RECT  2.370 0.465 2.480 3.440 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFCNQD2BWP7T

MACRO SDFD0BWP7T
    CLASS CORE ;
    FOREIGN SDFD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.075 13.300 2.560 ;
        RECT  12.885 1.075 13.020 1.305 ;
        RECT  12.600 2.330 13.020 2.560 ;
        RECT  12.655 0.520 12.885 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.510 14.420 2.715 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.470 1.760 4.620 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.660 0.810 ;
        RECT  10.530 -0.235 13.320 0.235 ;
        RECT  10.190 -0.235 10.530 0.465 ;
        RECT  8.510 -0.235 10.190 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.900 -0.235 4.575 0.235 ;
        RECT  3.560 -0.235 3.900 0.465 ;
        RECT  1.240 -0.235 3.560 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.730 3.685 14.560 4.155 ;
        RECT  13.390 3.365 13.730 4.155 ;
        RECT  11.430 3.685 13.390 4.155 ;
        RECT  11.090 3.385 11.430 4.155 ;
        RECT  8.520 3.685 11.090 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.960 3.685 8.160 4.155 ;
        RECT  4.620 3.455 4.960 4.155 ;
        RECT  3.780 3.685 4.620 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.240 3.685 3.440 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.020 ;
        RECT  12.370 2.790 13.615 3.020 ;
        RECT  10.990 0.465 12.420 0.695 ;
        RECT  12.140 1.020 12.370 3.020 ;
        RECT  11.450 1.020 12.140 1.250 ;
        RECT  11.900 2.540 12.140 2.775 ;
        RECT  11.680 1.565 11.910 2.310 ;
        RECT  11.450 2.080 11.680 2.310 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  11.220 2.080 11.450 2.995 ;
        RECT  10.735 1.600 11.220 1.830 ;
        RECT  9.935 2.765 11.220 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.500 2.300 10.770 2.530 ;
        RECT  10.500 0.990 10.760 1.220 ;
        RECT  10.270 0.990 10.500 2.530 ;
        RECT  9.225 3.225 10.480 3.455 ;
        RECT  9.705 0.910 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.375 ;
        RECT  5.845 3.145 7.520 3.375 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.615 6.080 1.955 ;
        RECT  5.615 0.925 5.845 3.375 ;
        RECT  5.375 2.560 5.615 2.790 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.090 ;
        RECT  2.600 0.695 5.145 0.925 ;
        RECT  4.240 1.155 5.140 1.385 ;
        RECT  4.240 2.505 4.345 2.845 ;
        RECT  4.010 1.155 4.240 2.845 ;
        RECT  2.445 0.695 2.600 2.780 ;
        RECT  2.370 0.695 2.445 3.355 ;
        RECT  2.195 0.695 2.370 0.925 ;
        RECT  2.215 2.545 2.370 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFD0BWP7T

MACRO SDFD1BWP7T
    CLASS CORE ;
    FOREIGN SDFD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.075 13.300 2.560 ;
        RECT  12.885 1.075 13.020 1.305 ;
        RECT  12.600 2.330 13.020 2.560 ;
        RECT  12.655 0.480 12.885 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.470 14.420 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.470 1.760 4.620 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.660 0.810 ;
        RECT  10.530 -0.235 13.320 0.235 ;
        RECT  10.190 -0.235 10.530 0.465 ;
        RECT  8.510 -0.235 10.190 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.900 -0.235 4.575 0.235 ;
        RECT  3.560 -0.235 3.900 0.465 ;
        RECT  1.240 -0.235 3.560 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 3.685 14.560 4.155 ;
        RECT  13.320 3.250 13.660 4.155 ;
        RECT  11.520 3.685 13.320 4.155 ;
        RECT  11.180 3.250 11.520 4.155 ;
        RECT  8.520 3.685 11.180 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.960 3.685 8.160 4.155 ;
        RECT  4.620 3.455 4.960 4.155 ;
        RECT  3.780 3.685 4.620 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.240 3.685 3.440 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.020 ;
        RECT  12.370 2.790 13.615 3.020 ;
        RECT  10.990 0.465 12.420 0.695 ;
        RECT  12.185 1.020 12.370 3.020 ;
        RECT  12.140 1.020 12.185 3.380 ;
        RECT  11.450 1.020 12.140 1.250 ;
        RECT  11.955 2.565 12.140 3.380 ;
        RECT  11.680 1.565 11.910 2.310 ;
        RECT  11.450 2.080 11.680 2.310 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  11.220 2.080 11.450 2.995 ;
        RECT  10.735 1.600 11.220 1.830 ;
        RECT  9.935 2.765 11.220 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.500 2.300 10.770 2.530 ;
        RECT  10.500 0.990 10.760 1.220 ;
        RECT  10.270 0.990 10.500 2.530 ;
        RECT  9.225 3.225 10.480 3.455 ;
        RECT  9.705 0.910 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.375 ;
        RECT  5.845 3.145 7.520 3.375 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.615 6.080 1.955 ;
        RECT  5.615 0.925 5.845 3.375 ;
        RECT  5.375 2.560 5.615 2.790 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.090 ;
        RECT  2.600 0.695 5.145 0.925 ;
        RECT  4.240 1.155 5.140 1.385 ;
        RECT  4.240 2.505 4.345 2.845 ;
        RECT  4.010 1.155 4.240 2.845 ;
        RECT  2.445 0.695 2.600 2.780 ;
        RECT  2.370 0.695 2.445 3.355 ;
        RECT  2.195 0.695 2.370 0.925 ;
        RECT  2.215 2.545 2.370 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFD1BWP7T

MACRO SDFD2BWP7T
    CLASS CORE ;
    FOREIGN SDFD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.560 0.465 13.905 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.055 15.540 2.690 ;
        RECT  15.260 0.465 15.285 3.310 ;
        RECT  15.050 0.465 15.260 1.285 ;
        RECT  15.055 2.460 15.260 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.470 1.760 4.620 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.245 ;
        RECT  14.620 -0.235 15.775 0.235 ;
        RECT  14.280 -0.235 14.620 1.180 ;
        RECT  13.140 -0.235 14.280 0.235 ;
        RECT  12.800 -0.235 13.140 0.465 ;
        RECT  11.510 -0.235 12.800 0.235 ;
        RECT  11.170 -0.235 11.510 0.465 ;
        RECT  8.495 -0.235 11.170 0.235 ;
        RECT  8.155 -0.235 8.495 0.730 ;
        RECT  4.905 -0.235 8.155 0.235 ;
        RECT  4.565 -0.235 4.905 0.465 ;
        RECT  3.900 -0.235 4.565 0.235 ;
        RECT  3.560 -0.235 3.900 0.465 ;
        RECT  1.240 -0.235 3.560 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.255 16.005 4.155 ;
        RECT  14.620 3.685 15.775 4.155 ;
        RECT  14.280 3.250 14.620 4.155 ;
        RECT  13.140 3.685 14.280 4.155 ;
        RECT  12.800 3.250 13.140 4.155 ;
        RECT  11.510 3.685 12.800 4.155 ;
        RECT  11.170 3.250 11.510 4.155 ;
        RECT  8.465 3.685 11.170 4.155 ;
        RECT  8.105 3.190 8.465 4.155 ;
        RECT  4.960 3.685 8.105 4.155 ;
        RECT  4.620 3.455 4.960 4.155 ;
        RECT  3.780 3.685 4.620 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.240 3.685 3.440 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.575 1.605 14.805 3.010 ;
        RECT  12.710 2.780 14.575 3.010 ;
        RECT  13.090 0.695 13.320 1.945 ;
        RECT  10.990 0.695 13.090 0.925 ;
        RECT  12.480 1.155 12.710 3.010 ;
        RECT  11.580 1.155 12.480 1.385 ;
        RECT  12.285 2.565 12.480 3.010 ;
        RECT  12.055 2.565 12.285 3.380 ;
        RECT  11.945 1.675 12.175 2.310 ;
        RECT  11.530 2.080 11.945 2.310 ;
        RECT  11.350 1.155 11.580 1.830 ;
        RECT  11.300 2.080 11.530 2.995 ;
        RECT  10.725 1.600 11.350 1.830 ;
        RECT  9.920 2.765 11.300 2.995 ;
        RECT  10.760 0.695 10.990 1.220 ;
        RECT  10.460 0.990 10.760 1.220 ;
        RECT  10.460 2.300 10.750 2.530 ;
        RECT  10.230 0.990 10.460 2.530 ;
        RECT  9.225 3.225 10.365 3.455 ;
        RECT  9.685 0.910 9.920 2.995 ;
        RECT  9.220 0.960 9.450 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  8.160 0.960 9.220 1.190 ;
        RECT  8.880 2.270 9.220 2.500 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.640 1.560 8.975 1.900 ;
        RECT  8.410 1.560 8.640 2.415 ;
        RECT  7.250 2.185 8.410 2.415 ;
        RECT  7.930 0.960 8.160 1.890 ;
        RECT  7.520 2.730 7.750 3.375 ;
        RECT  5.830 3.145 7.520 3.375 ;
        RECT  7.085 0.935 7.250 2.415 ;
        RECT  7.020 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.020 2.905 ;
        RECT  6.300 0.465 6.530 2.850 ;
        RECT  5.365 0.465 6.300 0.695 ;
        RECT  6.080 2.620 6.300 2.850 ;
        RECT  5.830 1.615 6.070 1.955 ;
        RECT  5.600 0.925 5.830 3.375 ;
        RECT  5.375 2.560 5.600 2.790 ;
        RECT  5.140 1.155 5.370 2.090 ;
        RECT  5.135 0.465 5.365 0.925 ;
        RECT  4.240 1.155 5.140 1.385 ;
        RECT  2.600 0.695 5.135 0.925 ;
        RECT  4.240 2.505 4.345 2.845 ;
        RECT  4.010 1.155 4.240 2.845 ;
        RECT  2.445 0.695 2.600 2.780 ;
        RECT  2.370 0.695 2.445 3.355 ;
        RECT  2.195 0.695 2.370 0.925 ;
        RECT  2.215 2.545 2.370 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFD2BWP7T

MACRO SDFKCND0BWP7T
    CLASS CORE ;
    FOREIGN SDFKCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.700 1.075 14.980 2.660 ;
        RECT  14.565 1.075 14.700 1.305 ;
        RECT  14.280 2.430 14.700 2.660 ;
        RECT  14.335 0.515 14.565 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.770 0.505 16.100 2.715 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.715 3.350 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.760 7.140 2.710 ;
        RECT  6.620 1.760 6.860 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.340 -0.235 16.240 0.235 ;
        RECT  15.000 -0.235 15.340 0.810 ;
        RECT  13.130 -0.235 15.000 0.235 ;
        RECT  12.790 -0.235 13.130 0.465 ;
        RECT  10.520 -0.235 12.790 0.235 ;
        RECT  10.180 -0.235 10.520 0.730 ;
        RECT  6.895 -0.235 10.180 0.235 ;
        RECT  6.555 -0.235 6.895 0.465 ;
        RECT  6.095 -0.235 6.555 0.235 ;
        RECT  5.685 -0.235 6.095 0.465 ;
        RECT  4.565 -0.235 5.685 0.235 ;
        RECT  4.225 -0.235 4.565 0.940 ;
        RECT  1.265 -0.235 4.225 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.255 3.685 16.240 4.155 ;
        RECT  14.915 3.455 15.255 4.155 ;
        RECT  13.160 3.685 14.915 4.155 ;
        RECT  12.820 3.455 13.160 4.155 ;
        RECT  10.530 3.685 12.820 4.155 ;
        RECT  10.170 3.190 10.530 4.155 ;
        RECT  7.110 3.685 10.170 4.155 ;
        RECT  6.770 3.455 7.110 4.155 ;
        RECT  6.045 3.685 6.770 4.155 ;
        RECT  5.705 3.455 6.045 4.155 ;
        RECT  4.060 3.685 5.705 4.155 ;
        RECT  3.680 3.455 4.060 4.155 ;
        RECT  1.265 3.685 3.680 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.295 1.600 15.525 3.215 ;
        RECT  13.100 2.985 15.295 3.215 ;
        RECT  14.050 1.605 14.470 1.945 ;
        RECT  13.820 0.950 14.050 2.755 ;
        RECT  12.890 0.950 13.820 1.180 ;
        RECT  13.580 2.520 13.820 2.755 ;
        RECT  13.330 1.565 13.560 2.290 ;
        RECT  13.100 2.060 13.330 2.290 ;
        RECT  12.870 2.060 13.100 3.215 ;
        RECT  12.660 0.950 12.890 1.830 ;
        RECT  11.945 2.060 12.870 2.290 ;
        RECT  11.235 3.225 12.390 3.455 ;
        RECT  11.715 0.910 11.945 2.860 ;
        RECT  11.255 0.960 11.485 2.500 ;
        RECT  10.205 0.960 11.255 1.190 ;
        RECT  10.940 2.270 11.255 2.500 ;
        RECT  11.005 2.730 11.235 3.455 ;
        RECT  9.830 2.730 11.005 2.960 ;
        RECT  10.710 1.560 10.985 1.900 ;
        RECT  10.480 1.560 10.710 2.415 ;
        RECT  9.275 2.185 10.480 2.415 ;
        RECT  9.975 0.960 10.205 1.890 ;
        RECT  9.600 2.730 9.830 3.375 ;
        RECT  8.055 3.145 9.600 3.375 ;
        RECT  9.235 0.935 9.275 2.415 ;
        RECT  9.005 0.935 9.235 2.905 ;
        RECT  8.610 0.995 8.755 2.840 ;
        RECT  8.525 0.520 8.610 2.840 ;
        RECT  8.270 0.520 8.525 1.220 ;
        RECT  8.285 2.420 8.525 2.840 ;
        RECT  7.345 0.520 8.270 0.750 ;
        RECT  8.055 1.615 8.230 1.955 ;
        RECT  8.030 1.615 8.055 3.375 ;
        RECT  7.825 0.980 8.030 3.375 ;
        RECT  7.800 0.980 7.825 2.760 ;
        RECT  7.570 0.980 7.800 1.210 ;
        RECT  7.525 2.530 7.800 2.760 ;
        RECT  7.345 2.995 7.575 3.455 ;
        RECT  7.120 0.520 7.345 0.925 ;
        RECT  6.555 2.995 7.345 3.225 ;
        RECT  5.225 0.695 7.120 0.925 ;
        RECT  6.325 2.560 6.555 3.225 ;
        RECT  6.305 1.155 6.540 1.385 ;
        RECT  6.305 2.560 6.325 2.790 ;
        RECT  6.075 1.155 6.305 2.790 ;
        RECT  5.515 1.620 5.745 3.225 ;
        RECT  2.660 2.995 5.515 3.225 ;
        RECT  4.995 0.495 5.225 2.765 ;
        RECT  3.810 2.450 4.560 2.680 ;
        RECT  3.580 0.685 3.810 2.680 ;
        RECT  2.890 0.685 3.580 0.915 ;
        RECT  2.895 2.450 3.580 2.680 ;
        RECT  2.430 0.850 2.660 3.225 ;
        RECT  2.125 0.850 2.430 1.080 ;
        RECT  2.130 2.440 2.430 2.680 ;
        RECT  1.940 1.310 2.180 2.080 ;
        RECT  0.465 1.310 1.940 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKCND0BWP7T

MACRO SDFKCND1BWP7T
    CLASS CORE ;
    FOREIGN SDFKCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.700 1.075 14.980 2.560 ;
        RECT  14.565 1.075 14.700 1.305 ;
        RECT  14.280 2.330 14.700 2.560 ;
        RECT  14.335 0.480 14.565 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.770 0.470 16.100 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.650 3.350 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.760 7.140 2.710 ;
        RECT  6.620 1.760 6.860 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.340 -0.235 16.240 0.235 ;
        RECT  15.000 -0.235 15.340 0.810 ;
        RECT  13.130 -0.235 15.000 0.235 ;
        RECT  12.790 -0.235 13.130 0.465 ;
        RECT  10.520 -0.235 12.790 0.235 ;
        RECT  10.180 -0.235 10.520 0.730 ;
        RECT  6.895 -0.235 10.180 0.235 ;
        RECT  6.555 -0.235 6.895 0.465 ;
        RECT  6.095 -0.235 6.555 0.235 ;
        RECT  5.685 -0.235 6.095 0.465 ;
        RECT  4.565 -0.235 5.685 0.235 ;
        RECT  4.225 -0.235 4.565 0.940 ;
        RECT  1.265 -0.235 4.225 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.340 3.685 16.240 4.155 ;
        RECT  15.000 3.250 15.340 4.155 ;
        RECT  13.160 3.685 15.000 4.155 ;
        RECT  12.820 3.455 13.160 4.155 ;
        RECT  10.530 3.685 12.820 4.155 ;
        RECT  10.170 3.190 10.530 4.155 ;
        RECT  7.110 3.685 10.170 4.155 ;
        RECT  6.770 3.455 7.110 4.155 ;
        RECT  6.045 3.685 6.770 4.155 ;
        RECT  5.705 3.455 6.045 4.155 ;
        RECT  4.060 3.685 5.705 4.155 ;
        RECT  3.680 3.455 4.060 4.155 ;
        RECT  1.265 3.685 3.680 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.295 1.600 15.525 3.020 ;
        RECT  14.665 2.790 15.295 3.020 ;
        RECT  14.435 2.790 14.665 3.215 ;
        RECT  14.050 1.605 14.470 1.945 ;
        RECT  13.100 2.985 14.435 3.215 ;
        RECT  13.820 0.950 14.050 2.755 ;
        RECT  12.890 0.950 13.820 1.180 ;
        RECT  13.580 2.520 13.820 2.755 ;
        RECT  13.330 1.565 13.560 2.290 ;
        RECT  13.100 2.060 13.330 2.290 ;
        RECT  12.870 2.060 13.100 3.215 ;
        RECT  12.660 0.950 12.890 1.825 ;
        RECT  11.945 2.060 12.870 2.290 ;
        RECT  11.235 3.225 12.390 3.455 ;
        RECT  11.715 0.910 11.945 2.860 ;
        RECT  11.255 0.960 11.485 2.500 ;
        RECT  10.205 0.960 11.255 1.190 ;
        RECT  10.940 2.270 11.255 2.500 ;
        RECT  11.005 2.730 11.235 3.455 ;
        RECT  9.830 2.730 11.005 2.960 ;
        RECT  10.710 1.560 10.985 1.900 ;
        RECT  10.480 1.560 10.710 2.415 ;
        RECT  9.275 2.185 10.480 2.415 ;
        RECT  9.975 0.960 10.205 1.890 ;
        RECT  9.600 2.730 9.830 3.375 ;
        RECT  8.055 3.145 9.600 3.375 ;
        RECT  9.235 0.935 9.275 2.415 ;
        RECT  9.005 0.935 9.235 2.905 ;
        RECT  8.610 1.005 8.755 2.840 ;
        RECT  8.525 0.520 8.610 2.840 ;
        RECT  8.270 0.520 8.525 1.220 ;
        RECT  8.285 2.420 8.525 2.840 ;
        RECT  7.345 0.520 8.270 0.750 ;
        RECT  8.055 1.615 8.230 1.955 ;
        RECT  8.030 1.615 8.055 3.375 ;
        RECT  7.825 0.980 8.030 3.375 ;
        RECT  7.800 0.980 7.825 2.760 ;
        RECT  7.570 0.980 7.800 1.210 ;
        RECT  7.525 2.530 7.800 2.760 ;
        RECT  7.345 2.995 7.575 3.455 ;
        RECT  7.120 0.520 7.345 0.925 ;
        RECT  6.555 2.995 7.345 3.225 ;
        RECT  5.225 0.695 7.120 0.925 ;
        RECT  6.325 2.560 6.555 3.225 ;
        RECT  6.305 1.155 6.540 1.385 ;
        RECT  6.305 2.560 6.325 2.790 ;
        RECT  6.075 1.155 6.305 2.790 ;
        RECT  5.515 1.620 5.745 3.225 ;
        RECT  2.660 2.995 5.515 3.225 ;
        RECT  4.995 0.495 5.225 2.765 ;
        RECT  3.810 2.450 4.560 2.680 ;
        RECT  3.580 0.685 3.810 2.680 ;
        RECT  2.890 0.685 3.580 0.915 ;
        RECT  2.895 2.450 3.580 2.680 ;
        RECT  2.430 0.850 2.660 3.225 ;
        RECT  2.125 0.850 2.430 1.080 ;
        RECT  2.130 2.440 2.430 2.680 ;
        RECT  1.940 1.310 2.180 2.080 ;
        RECT  0.465 1.310 1.940 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKCND1BWP7T

MACRO SDFKCND2BWP7T
    CLASS CORE ;
    FOREIGN SDFKCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3346 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.240 0.490 15.580 2.560 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 1.060 17.220 2.735 ;
        RECT  16.940 0.480 16.965 3.310 ;
        RECT  16.735 0.480 16.940 1.290 ;
        RECT  16.735 2.500 16.940 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.715 3.350 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.760 7.140 2.710 ;
        RECT  6.620 1.760 6.860 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 -0.235 17.920 0.235 ;
        RECT  17.455 -0.235 17.685 1.275 ;
        RECT  16.300 -0.235 17.455 0.235 ;
        RECT  15.960 -0.235 16.300 1.190 ;
        RECT  14.820 -0.235 15.960 0.235 ;
        RECT  14.480 -0.235 14.820 1.190 ;
        RECT  13.355 -0.235 14.480 0.235 ;
        RECT  13.015 -0.235 13.355 0.670 ;
        RECT  10.520 -0.235 13.015 0.235 ;
        RECT  10.180 -0.235 10.520 0.730 ;
        RECT  6.895 -0.235 10.180 0.235 ;
        RECT  6.555 -0.235 6.895 0.465 ;
        RECT  6.095 -0.235 6.555 0.235 ;
        RECT  5.685 -0.235 6.095 0.465 ;
        RECT  4.565 -0.235 5.685 0.235 ;
        RECT  4.225 -0.235 4.565 0.940 ;
        RECT  1.265 -0.235 4.225 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 3.685 17.920 4.155 ;
        RECT  17.455 2.255 17.685 4.155 ;
        RECT  16.300 3.685 17.455 4.155 ;
        RECT  15.960 3.250 16.300 4.155 ;
        RECT  14.740 3.685 15.960 4.155 ;
        RECT  14.400 3.455 14.740 4.155 ;
        RECT  13.225 3.685 14.400 4.155 ;
        RECT  12.885 3.455 13.225 4.155 ;
        RECT  10.530 3.685 12.885 4.155 ;
        RECT  10.170 3.190 10.530 4.155 ;
        RECT  7.110 3.685 10.170 4.155 ;
        RECT  6.770 3.455 7.110 4.155 ;
        RECT  6.045 3.685 6.770 4.155 ;
        RECT  5.705 3.455 6.045 4.155 ;
        RECT  4.060 3.685 5.705 4.155 ;
        RECT  3.680 3.455 4.060 4.155 ;
        RECT  1.265 3.685 3.680 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.255 1.600 16.485 3.020 ;
        RECT  14.950 2.790 16.255 3.020 ;
        RECT  14.040 1.615 15.010 1.955 ;
        RECT  14.720 2.790 14.950 3.215 ;
        RECT  13.100 2.985 14.720 3.215 ;
        RECT  13.810 0.465 14.040 2.755 ;
        RECT  12.890 0.940 13.810 1.170 ;
        RECT  13.690 2.520 13.810 2.755 ;
        RECT  13.330 1.565 13.560 2.290 ;
        RECT  13.100 2.060 13.330 2.290 ;
        RECT  12.870 2.060 13.100 3.215 ;
        RECT  12.660 0.940 12.890 1.830 ;
        RECT  11.945 2.060 12.870 2.290 ;
        RECT  11.235 3.225 12.390 3.455 ;
        RECT  11.715 0.910 11.945 2.860 ;
        RECT  11.235 0.960 11.465 2.500 ;
        RECT  10.205 0.960 11.235 1.190 ;
        RECT  10.940 2.270 11.235 2.500 ;
        RECT  11.005 2.730 11.235 3.455 ;
        RECT  9.830 2.730 11.005 2.960 ;
        RECT  10.710 1.560 10.985 1.900 ;
        RECT  10.480 1.560 10.710 2.415 ;
        RECT  9.275 2.185 10.480 2.415 ;
        RECT  9.975 0.960 10.205 1.890 ;
        RECT  9.600 2.730 9.830 3.375 ;
        RECT  8.055 3.145 9.600 3.375 ;
        RECT  9.235 0.935 9.275 2.415 ;
        RECT  9.005 0.935 9.235 2.905 ;
        RECT  8.610 1.000 8.755 2.840 ;
        RECT  8.525 0.520 8.610 2.840 ;
        RECT  8.270 0.520 8.525 1.220 ;
        RECT  8.285 2.420 8.525 2.840 ;
        RECT  7.345 0.520 8.270 0.750 ;
        RECT  8.055 1.615 8.230 1.955 ;
        RECT  8.030 1.615 8.055 3.375 ;
        RECT  7.825 0.980 8.030 3.375 ;
        RECT  7.800 0.980 7.825 2.760 ;
        RECT  7.570 0.980 7.800 1.210 ;
        RECT  7.525 2.530 7.800 2.760 ;
        RECT  7.345 2.995 7.575 3.455 ;
        RECT  7.120 0.520 7.345 0.925 ;
        RECT  6.555 2.995 7.345 3.225 ;
        RECT  5.225 0.695 7.120 0.925 ;
        RECT  6.325 2.560 6.555 3.225 ;
        RECT  6.305 1.155 6.540 1.385 ;
        RECT  6.305 2.560 6.325 2.790 ;
        RECT  6.075 1.155 6.305 2.790 ;
        RECT  5.515 1.620 5.745 3.225 ;
        RECT  2.660 2.995 5.515 3.225 ;
        RECT  4.995 0.495 5.225 2.765 ;
        RECT  3.810 2.450 4.560 2.680 ;
        RECT  3.580 0.685 3.810 2.680 ;
        RECT  2.890 0.685 3.580 0.915 ;
        RECT  2.895 2.450 3.580 2.680 ;
        RECT  2.430 0.850 2.660 3.225 ;
        RECT  2.125 0.850 2.430 1.080 ;
        RECT  2.130 2.440 2.430 2.680 ;
        RECT  1.940 1.310 2.180 2.080 ;
        RECT  0.465 1.310 1.940 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKCND2BWP7T

MACRO SDFKCNQD0BWP7T
    CLASS CORE ;
    FOREIGN SDFKCNQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.210 0.640 15.540 2.965 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.715 3.350 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.760 7.140 2.710 ;
        RECT  6.620 1.760 6.860 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.725 -0.235 15.680 0.235 ;
        RECT  14.495 -0.235 14.725 0.990 ;
        RECT  13.300 -0.235 14.495 0.235 ;
        RECT  12.960 -0.235 13.300 0.720 ;
        RECT  10.520 -0.235 12.960 0.235 ;
        RECT  10.180 -0.235 10.520 0.730 ;
        RECT  6.895 -0.235 10.180 0.235 ;
        RECT  6.555 -0.235 6.895 0.465 ;
        RECT  6.095 -0.235 6.555 0.235 ;
        RECT  5.685 -0.235 6.095 0.465 ;
        RECT  4.565 -0.235 5.685 0.235 ;
        RECT  4.225 -0.235 4.565 0.940 ;
        RECT  1.265 -0.235 4.225 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.725 3.685 15.680 4.155 ;
        RECT  14.495 2.615 14.725 4.155 ;
        RECT  13.320 3.685 14.495 4.155 ;
        RECT  12.980 2.665 13.320 4.155 ;
        RECT  10.530 3.685 12.980 4.155 ;
        RECT  10.170 3.190 10.530 4.155 ;
        RECT  7.110 3.685 10.170 4.155 ;
        RECT  6.770 3.455 7.110 4.155 ;
        RECT  6.045 3.685 6.770 4.155 ;
        RECT  5.705 3.455 6.045 4.155 ;
        RECT  4.060 3.685 5.705 4.155 ;
        RECT  3.680 3.455 4.060 4.155 ;
        RECT  1.265 3.685 3.680 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.030 0.950 14.260 2.915 ;
        RECT  12.890 0.950 14.030 1.180 ;
        RECT  13.740 2.680 14.030 2.915 ;
        RECT  13.555 1.660 13.785 2.360 ;
        RECT  11.945 2.130 13.555 2.360 ;
        RECT  12.660 0.950 12.890 1.830 ;
        RECT  11.235 3.225 12.370 3.455 ;
        RECT  11.715 0.910 11.945 2.850 ;
        RECT  11.255 0.960 11.485 2.500 ;
        RECT  10.205 0.960 11.255 1.190 ;
        RECT  10.940 2.270 11.255 2.500 ;
        RECT  11.005 2.730 11.235 3.455 ;
        RECT  9.830 2.730 11.005 2.960 ;
        RECT  10.710 1.560 10.985 1.900 ;
        RECT  10.480 1.560 10.710 2.415 ;
        RECT  9.275 2.185 10.480 2.415 ;
        RECT  9.975 0.960 10.205 1.890 ;
        RECT  9.600 2.730 9.830 3.375 ;
        RECT  8.055 3.145 9.600 3.375 ;
        RECT  9.235 0.935 9.275 2.415 ;
        RECT  9.005 0.935 9.235 2.905 ;
        RECT  8.610 1.000 8.755 2.840 ;
        RECT  8.525 0.520 8.610 2.840 ;
        RECT  8.270 0.520 8.525 1.220 ;
        RECT  8.285 2.420 8.525 2.840 ;
        RECT  7.345 0.520 8.270 0.750 ;
        RECT  8.055 1.615 8.230 1.955 ;
        RECT  8.030 1.615 8.055 3.375 ;
        RECT  7.825 0.980 8.030 3.375 ;
        RECT  7.800 0.980 7.825 2.760 ;
        RECT  7.570 0.980 7.800 1.210 ;
        RECT  7.525 2.530 7.800 2.760 ;
        RECT  7.345 2.995 7.575 3.455 ;
        RECT  7.120 0.520 7.345 0.925 ;
        RECT  6.555 2.995 7.345 3.225 ;
        RECT  5.225 0.695 7.120 0.925 ;
        RECT  6.325 2.560 6.555 3.225 ;
        RECT  6.305 1.155 6.540 1.385 ;
        RECT  6.305 2.560 6.325 2.790 ;
        RECT  6.075 1.155 6.305 2.790 ;
        RECT  5.515 1.620 5.745 3.225 ;
        RECT  2.660 2.995 5.515 3.225 ;
        RECT  4.995 0.495 5.225 2.765 ;
        RECT  3.810 2.450 4.560 2.680 ;
        RECT  3.580 0.685 3.810 2.680 ;
        RECT  2.890 0.685 3.580 0.915 ;
        RECT  2.895 2.450 3.580 2.680 ;
        RECT  2.430 0.850 2.660 3.225 ;
        RECT  2.125 0.850 2.430 1.080 ;
        RECT  2.130 2.440 2.430 2.680 ;
        RECT  1.940 1.310 2.180 2.080 ;
        RECT  0.465 1.310 1.940 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKCNQD0BWP7T

MACRO SDFKCNQD1BWP7T
    CLASS CORE ;
    FOREIGN SDFKCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.210 0.470 15.540 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.715 3.350 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.760 7.140 2.710 ;
        RECT  6.620 1.760 6.860 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.725 -0.235 15.680 0.235 ;
        RECT  14.495 -0.235 14.725 1.245 ;
        RECT  13.300 -0.235 14.495 0.235 ;
        RECT  12.960 -0.235 13.300 0.720 ;
        RECT  10.520 -0.235 12.960 0.235 ;
        RECT  10.180 -0.235 10.520 0.730 ;
        RECT  6.895 -0.235 10.180 0.235 ;
        RECT  6.555 -0.235 6.895 0.465 ;
        RECT  6.095 -0.235 6.555 0.235 ;
        RECT  5.685 -0.235 6.095 0.465 ;
        RECT  4.565 -0.235 5.685 0.235 ;
        RECT  4.225 -0.235 4.565 0.940 ;
        RECT  1.265 -0.235 4.225 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.725 3.685 15.680 4.155 ;
        RECT  14.495 2.255 14.725 4.155 ;
        RECT  13.320 3.685 14.495 4.155 ;
        RECT  12.980 2.665 13.320 4.155 ;
        RECT  10.530 3.685 12.980 4.155 ;
        RECT  10.170 3.190 10.530 4.155 ;
        RECT  7.110 3.685 10.170 4.155 ;
        RECT  6.770 3.455 7.110 4.155 ;
        RECT  6.045 3.685 6.770 4.155 ;
        RECT  5.705 3.455 6.045 4.155 ;
        RECT  4.060 3.685 5.705 4.155 ;
        RECT  3.680 3.455 4.060 4.155 ;
        RECT  1.265 3.685 3.680 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.035 0.950 14.265 2.915 ;
        RECT  12.890 0.950 14.035 1.180 ;
        RECT  13.740 2.680 14.035 2.915 ;
        RECT  13.555 1.600 13.785 2.290 ;
        RECT  11.945 2.060 13.555 2.290 ;
        RECT  12.660 0.950 12.890 1.830 ;
        RECT  11.235 3.225 12.370 3.455 ;
        RECT  11.715 0.910 11.945 2.850 ;
        RECT  11.255 0.960 11.485 2.500 ;
        RECT  10.205 0.960 11.255 1.190 ;
        RECT  10.940 2.270 11.255 2.500 ;
        RECT  11.005 2.730 11.235 3.455 ;
        RECT  9.830 2.730 11.005 2.960 ;
        RECT  10.710 1.560 10.985 1.900 ;
        RECT  10.480 1.560 10.710 2.415 ;
        RECT  9.275 2.185 10.480 2.415 ;
        RECT  9.975 0.960 10.205 1.890 ;
        RECT  9.600 2.730 9.830 3.375 ;
        RECT  8.055 3.145 9.600 3.375 ;
        RECT  9.235 0.935 9.275 2.415 ;
        RECT  9.005 0.935 9.235 2.905 ;
        RECT  8.610 1.005 8.755 2.840 ;
        RECT  8.525 0.520 8.610 2.840 ;
        RECT  8.270 0.520 8.525 1.220 ;
        RECT  8.285 2.420 8.525 2.840 ;
        RECT  7.345 0.520 8.270 0.750 ;
        RECT  8.055 1.615 8.230 1.955 ;
        RECT  8.030 1.615 8.055 3.375 ;
        RECT  7.825 0.980 8.030 3.375 ;
        RECT  7.800 0.980 7.825 2.760 ;
        RECT  7.570 0.980 7.800 1.210 ;
        RECT  7.525 2.530 7.800 2.760 ;
        RECT  7.345 2.995 7.575 3.455 ;
        RECT  7.120 0.520 7.345 0.925 ;
        RECT  6.555 2.995 7.345 3.225 ;
        RECT  5.225 0.695 7.120 0.925 ;
        RECT  6.325 2.560 6.555 3.225 ;
        RECT  6.305 1.155 6.540 1.385 ;
        RECT  6.305 2.560 6.325 2.790 ;
        RECT  6.075 1.155 6.305 2.790 ;
        RECT  5.515 1.620 5.745 3.225 ;
        RECT  2.660 2.995 5.515 3.225 ;
        RECT  4.995 0.495 5.225 2.765 ;
        RECT  3.810 2.450 4.560 2.680 ;
        RECT  3.580 0.685 3.810 2.680 ;
        RECT  2.890 0.685 3.580 0.915 ;
        RECT  2.895 2.450 3.580 2.680 ;
        RECT  2.430 0.850 2.660 3.225 ;
        RECT  2.125 0.850 2.430 1.080 ;
        RECT  2.130 2.440 2.430 2.680 ;
        RECT  1.940 1.310 2.180 2.080 ;
        RECT  0.465 1.310 1.940 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKCNQD1BWP7T

MACRO SDFKCNQD2BWP7T
    CLASS CORE ;
    FOREIGN SDFKCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.060 15.540 2.725 ;
        RECT  15.260 0.470 15.285 3.310 ;
        RECT  15.055 0.470 15.260 1.290 ;
        RECT  15.055 2.495 15.260 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.715 3.350 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.860 1.760 7.140 2.710 ;
        RECT  6.620 1.760 6.860 2.105 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.2556 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.245 ;
        RECT  14.565 -0.235 15.775 0.235 ;
        RECT  14.335 -0.235 14.565 1.245 ;
        RECT  13.125 -0.235 14.335 0.235 ;
        RECT  12.785 -0.235 13.125 0.465 ;
        RECT  10.520 -0.235 12.785 0.235 ;
        RECT  10.180 -0.235 10.520 0.730 ;
        RECT  6.895 -0.235 10.180 0.235 ;
        RECT  6.555 -0.235 6.895 0.465 ;
        RECT  6.095 -0.235 6.555 0.235 ;
        RECT  5.685 -0.235 6.095 0.465 ;
        RECT  4.565 -0.235 5.685 0.235 ;
        RECT  4.225 -0.235 4.565 0.940 ;
        RECT  1.265 -0.235 4.225 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.255 16.005 4.155 ;
        RECT  14.565 3.685 15.775 4.155 ;
        RECT  14.335 2.255 14.565 4.155 ;
        RECT  13.135 3.685 14.335 4.155 ;
        RECT  12.795 3.350 13.135 4.155 ;
        RECT  10.530 3.685 12.795 4.155 ;
        RECT  10.170 3.190 10.530 4.155 ;
        RECT  7.110 3.685 10.170 4.155 ;
        RECT  6.770 3.455 7.110 4.155 ;
        RECT  6.045 3.685 6.770 4.155 ;
        RECT  5.705 3.455 6.045 4.155 ;
        RECT  4.060 3.685 5.705 4.155 ;
        RECT  3.680 3.455 4.060 4.155 ;
        RECT  1.265 3.685 3.680 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.875 0.950 14.105 2.915 ;
        RECT  12.890 0.950 13.875 1.180 ;
        RECT  13.580 2.680 13.875 2.915 ;
        RECT  13.395 1.610 13.625 2.410 ;
        RECT  11.945 2.180 13.395 2.410 ;
        RECT  12.660 0.950 12.890 1.905 ;
        RECT  11.235 3.225 12.370 3.455 ;
        RECT  11.715 0.910 11.945 2.850 ;
        RECT  11.255 0.960 11.485 2.500 ;
        RECT  10.205 0.960 11.255 1.190 ;
        RECT  10.940 2.270 11.255 2.500 ;
        RECT  11.005 2.730 11.235 3.455 ;
        RECT  9.830 2.730 11.005 2.960 ;
        RECT  10.710 1.560 10.985 1.900 ;
        RECT  10.480 1.560 10.710 2.415 ;
        RECT  9.275 2.185 10.480 2.415 ;
        RECT  9.975 0.960 10.205 1.890 ;
        RECT  9.600 2.730 9.830 3.375 ;
        RECT  8.055 3.145 9.600 3.375 ;
        RECT  9.235 0.935 9.275 2.415 ;
        RECT  9.005 0.935 9.235 2.905 ;
        RECT  8.610 1.005 8.755 2.840 ;
        RECT  8.525 0.520 8.610 2.840 ;
        RECT  8.270 0.520 8.525 1.220 ;
        RECT  8.285 2.420 8.525 2.840 ;
        RECT  7.345 0.520 8.270 0.750 ;
        RECT  8.055 1.615 8.230 1.955 ;
        RECT  8.030 1.615 8.055 3.375 ;
        RECT  7.825 0.980 8.030 3.375 ;
        RECT  7.800 0.980 7.825 2.760 ;
        RECT  7.570 0.980 7.800 1.210 ;
        RECT  7.525 2.530 7.800 2.760 ;
        RECT  7.345 2.995 7.575 3.455 ;
        RECT  7.120 0.520 7.345 0.925 ;
        RECT  6.555 2.995 7.345 3.225 ;
        RECT  5.225 0.695 7.120 0.925 ;
        RECT  6.325 2.560 6.555 3.225 ;
        RECT  6.305 1.155 6.540 1.385 ;
        RECT  6.305 2.560 6.325 2.790 ;
        RECT  6.075 1.155 6.305 2.790 ;
        RECT  5.515 1.620 5.745 3.225 ;
        RECT  2.660 2.995 5.515 3.225 ;
        RECT  4.995 0.495 5.225 2.765 ;
        RECT  3.810 2.450 4.560 2.680 ;
        RECT  3.580 0.685 3.810 2.680 ;
        RECT  2.890 0.685 3.580 0.915 ;
        RECT  2.895 2.450 3.580 2.680 ;
        RECT  2.430 0.850 2.660 3.225 ;
        RECT  2.125 0.850 2.430 1.080 ;
        RECT  2.130 2.440 2.430 2.680 ;
        RECT  1.940 1.310 2.180 2.080 ;
        RECT  0.465 1.310 1.940 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKCNQD2BWP7T

MACRO SDFKSND0BWP7T
    CLASS CORE ;
    FOREIGN SDFKSND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.210 5.460 2.150 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.820 1.075 16.100 2.645 ;
        RECT  15.685 1.075 15.820 1.305 ;
        RECT  15.400 2.415 15.820 2.645 ;
        RECT  15.455 0.480 15.685 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.890 0.470 17.220 2.715 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.680 3.420 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.760 8.260 2.710 ;
        RECT  7.740 1.760 7.980 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.460 -0.235 17.360 0.235 ;
        RECT  16.120 -0.235 16.460 0.775 ;
        RECT  14.220 -0.235 16.120 0.235 ;
        RECT  13.880 -0.235 14.220 0.465 ;
        RECT  11.640 -0.235 13.880 0.235 ;
        RECT  11.300 -0.235 11.640 0.730 ;
        RECT  8.015 -0.235 11.300 0.235 ;
        RECT  7.675 -0.235 8.015 0.465 ;
        RECT  7.225 -0.235 7.675 0.235 ;
        RECT  6.815 -0.235 7.225 0.465 ;
        RECT  3.945 -0.235 6.815 0.235 ;
        RECT  3.605 -0.235 3.945 0.465 ;
        RECT  1.265 -0.235 3.605 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.395 3.685 17.360 4.155 ;
        RECT  16.055 3.455 16.395 4.155 ;
        RECT  14.280 3.685 16.055 4.155 ;
        RECT  13.940 3.455 14.280 4.155 ;
        RECT  11.650 3.685 13.940 4.155 ;
        RECT  11.290 3.190 11.650 4.155 ;
        RECT  8.230 3.685 11.290 4.155 ;
        RECT  7.890 3.455 8.230 4.155 ;
        RECT  7.170 3.685 7.890 4.155 ;
        RECT  6.830 3.455 7.170 4.155 ;
        RECT  4.775 3.685 6.830 4.155 ;
        RECT  4.435 3.455 4.775 4.155 ;
        RECT  1.265 3.685 4.435 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.415 1.600 16.645 3.215 ;
        RECT  14.220 2.985 16.415 3.215 ;
        RECT  15.170 1.605 15.590 1.945 ;
        RECT  14.940 0.950 15.170 2.750 ;
        RECT  14.010 0.950 14.940 1.180 ;
        RECT  14.700 2.520 14.940 2.750 ;
        RECT  14.450 1.515 14.680 2.290 ;
        RECT  14.220 2.060 14.450 2.290 ;
        RECT  13.990 2.060 14.220 3.215 ;
        RECT  13.780 0.950 14.010 1.830 ;
        RECT  13.065 2.060 13.990 2.290 ;
        RECT  12.355 3.225 13.510 3.455 ;
        RECT  12.835 0.910 13.065 2.860 ;
        RECT  12.375 0.960 12.605 2.500 ;
        RECT  11.325 0.960 12.375 1.190 ;
        RECT  12.060 2.270 12.375 2.500 ;
        RECT  12.125 2.730 12.355 3.455 ;
        RECT  10.950 2.730 12.125 2.960 ;
        RECT  11.830 1.560 12.105 1.900 ;
        RECT  11.600 1.560 11.830 2.415 ;
        RECT  10.395 2.185 11.600 2.415 ;
        RECT  11.095 0.960 11.325 1.890 ;
        RECT  10.720 2.730 10.950 3.375 ;
        RECT  9.175 3.145 10.720 3.375 ;
        RECT  10.355 0.935 10.395 2.415 ;
        RECT  10.125 0.935 10.355 2.905 ;
        RECT  9.730 0.990 9.875 2.840 ;
        RECT  9.645 0.520 9.730 2.840 ;
        RECT  9.390 0.520 9.645 1.220 ;
        RECT  9.405 2.420 9.645 2.840 ;
        RECT  8.465 0.520 9.390 0.750 ;
        RECT  9.175 1.615 9.350 1.955 ;
        RECT  9.150 1.615 9.175 3.375 ;
        RECT  8.945 0.980 9.150 3.375 ;
        RECT  8.920 0.980 8.945 2.760 ;
        RECT  8.690 0.980 8.920 1.210 ;
        RECT  8.645 2.530 8.920 2.760 ;
        RECT  8.465 2.995 8.695 3.455 ;
        RECT  8.240 0.520 8.465 0.925 ;
        RECT  7.675 2.995 8.465 3.225 ;
        RECT  6.355 0.695 8.240 0.925 ;
        RECT  7.445 2.560 7.675 3.225 ;
        RECT  7.425 1.155 7.670 1.385 ;
        RECT  7.425 2.560 7.445 2.790 ;
        RECT  7.195 1.155 7.425 2.790 ;
        RECT  6.645 1.620 6.875 3.225 ;
        RECT  2.615 2.995 6.645 3.225 ;
        RECT  6.115 0.495 6.355 2.765 ;
        RECT  4.870 0.480 5.710 0.710 ;
        RECT  4.870 2.450 5.680 2.680 ;
        RECT  4.640 0.480 4.870 2.680 ;
        RECT  4.185 1.665 4.640 1.895 ;
        RECT  3.930 1.020 4.390 1.250 ;
        RECT  3.700 0.750 3.930 2.680 ;
        RECT  3.075 0.750 3.700 0.980 ;
        RECT  2.940 2.450 3.700 2.680 ;
        RECT  2.845 0.510 3.075 0.980 ;
        RECT  2.385 0.850 2.615 3.225 ;
        RECT  2.050 0.850 2.385 1.080 ;
        RECT  2.130 2.440 2.385 2.680 ;
        RECT  1.925 1.310 2.155 2.080 ;
        RECT  0.465 1.310 1.925 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKSND0BWP7T

MACRO SDFKSND1BWP7T
    CLASS CORE ;
    FOREIGN SDFKSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.210 5.460 2.150 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.820 1.075 16.100 2.560 ;
        RECT  15.685 1.075 15.820 1.305 ;
        RECT  15.400 2.330 15.820 2.560 ;
        RECT  15.455 0.480 15.685 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.890 0.470 17.220 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.680 3.420 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.760 8.260 2.710 ;
        RECT  7.740 1.760 7.980 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.460 -0.235 17.360 0.235 ;
        RECT  16.120 -0.235 16.460 0.810 ;
        RECT  14.235 -0.235 16.120 0.235 ;
        RECT  13.895 -0.235 14.235 0.465 ;
        RECT  11.640 -0.235 13.895 0.235 ;
        RECT  11.300 -0.235 11.640 0.730 ;
        RECT  8.015 -0.235 11.300 0.235 ;
        RECT  7.675 -0.235 8.015 0.465 ;
        RECT  7.225 -0.235 7.675 0.235 ;
        RECT  6.815 -0.235 7.225 0.465 ;
        RECT  3.945 -0.235 6.815 0.235 ;
        RECT  3.605 -0.235 3.945 0.465 ;
        RECT  1.265 -0.235 3.605 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.460 3.685 17.360 4.155 ;
        RECT  16.120 3.250 16.460 4.155 ;
        RECT  14.280 3.685 16.120 4.155 ;
        RECT  13.940 3.455 14.280 4.155 ;
        RECT  11.650 3.685 13.940 4.155 ;
        RECT  11.290 3.190 11.650 4.155 ;
        RECT  8.230 3.685 11.290 4.155 ;
        RECT  7.890 3.455 8.230 4.155 ;
        RECT  7.170 3.685 7.890 4.155 ;
        RECT  6.830 3.455 7.170 4.155 ;
        RECT  4.775 3.685 6.830 4.155 ;
        RECT  4.435 3.455 4.775 4.155 ;
        RECT  1.265 3.685 4.435 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.415 1.600 16.645 3.020 ;
        RECT  15.785 2.790 16.415 3.020 ;
        RECT  15.555 2.790 15.785 3.215 ;
        RECT  15.170 1.605 15.590 1.945 ;
        RECT  14.220 2.985 15.555 3.215 ;
        RECT  14.940 0.950 15.170 2.750 ;
        RECT  14.010 0.950 14.940 1.180 ;
        RECT  14.700 2.520 14.940 2.750 ;
        RECT  14.450 1.565 14.680 2.290 ;
        RECT  14.220 2.060 14.450 2.290 ;
        RECT  13.990 2.060 14.220 3.215 ;
        RECT  13.780 0.950 14.010 1.830 ;
        RECT  13.065 2.060 13.990 2.290 ;
        RECT  12.355 3.225 13.510 3.455 ;
        RECT  12.835 0.910 13.065 2.850 ;
        RECT  12.375 0.960 12.605 2.500 ;
        RECT  11.325 0.960 12.375 1.190 ;
        RECT  12.060 2.270 12.375 2.500 ;
        RECT  12.125 2.730 12.355 3.455 ;
        RECT  10.950 2.730 12.125 2.960 ;
        RECT  11.830 1.560 12.105 1.900 ;
        RECT  11.600 1.560 11.830 2.415 ;
        RECT  10.395 2.185 11.600 2.415 ;
        RECT  11.095 0.960 11.325 1.890 ;
        RECT  10.720 2.730 10.950 3.375 ;
        RECT  9.175 3.145 10.720 3.375 ;
        RECT  10.355 0.935 10.395 2.415 ;
        RECT  10.125 0.935 10.355 2.905 ;
        RECT  9.735 0.995 9.875 2.840 ;
        RECT  9.645 0.520 9.735 2.840 ;
        RECT  9.390 0.520 9.645 1.220 ;
        RECT  9.405 2.420 9.645 2.840 ;
        RECT  8.465 0.520 9.390 0.750 ;
        RECT  9.175 1.615 9.350 1.955 ;
        RECT  9.150 1.615 9.175 3.375 ;
        RECT  8.945 0.980 9.150 3.375 ;
        RECT  8.920 0.980 8.945 2.760 ;
        RECT  8.690 0.980 8.920 1.210 ;
        RECT  8.645 2.530 8.920 2.760 ;
        RECT  8.465 2.995 8.695 3.455 ;
        RECT  8.240 0.520 8.465 0.925 ;
        RECT  7.675 2.995 8.465 3.225 ;
        RECT  6.355 0.695 8.240 0.925 ;
        RECT  7.445 2.560 7.675 3.225 ;
        RECT  7.425 1.155 7.670 1.385 ;
        RECT  7.425 2.560 7.445 2.790 ;
        RECT  7.195 1.155 7.425 2.790 ;
        RECT  6.645 1.620 6.875 3.225 ;
        RECT  2.615 2.995 6.645 3.225 ;
        RECT  6.115 0.495 6.355 2.765 ;
        RECT  4.870 0.480 5.710 0.710 ;
        RECT  4.870 2.450 5.680 2.680 ;
        RECT  4.640 0.480 4.870 2.680 ;
        RECT  4.185 1.665 4.640 1.895 ;
        RECT  3.930 1.020 4.390 1.250 ;
        RECT  3.700 0.750 3.930 2.680 ;
        RECT  3.075 0.750 3.700 0.980 ;
        RECT  2.940 2.450 3.700 2.680 ;
        RECT  2.845 0.510 3.075 0.980 ;
        RECT  2.385 0.850 2.615 3.225 ;
        RECT  2.050 0.850 2.385 1.080 ;
        RECT  2.130 2.440 2.385 2.680 ;
        RECT  1.925 1.310 2.155 2.080 ;
        RECT  0.465 1.310 1.925 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKSND1BWP7T

MACRO SDFKSND2BWP7T
    CLASS CORE ;
    FOREIGN SDFKSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.210 5.460 2.150 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3346 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.360 0.490 16.700 2.560 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.085 1.060 18.340 2.735 ;
        RECT  18.060 0.480 18.085 3.310 ;
        RECT  17.855 0.480 18.060 1.290 ;
        RECT  17.855 2.500 18.060 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.680 3.420 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.760 8.260 2.710 ;
        RECT  7.740 1.760 7.980 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.805 -0.235 19.040 0.235 ;
        RECT  18.575 -0.235 18.805 1.275 ;
        RECT  17.420 -0.235 18.575 0.235 ;
        RECT  17.080 -0.235 17.420 1.190 ;
        RECT  15.940 -0.235 17.080 0.235 ;
        RECT  15.600 -0.235 15.940 1.190 ;
        RECT  14.475 -0.235 15.600 0.235 ;
        RECT  14.135 -0.235 14.475 0.670 ;
        RECT  11.640 -0.235 14.135 0.235 ;
        RECT  11.300 -0.235 11.640 0.730 ;
        RECT  8.015 -0.235 11.300 0.235 ;
        RECT  7.675 -0.235 8.015 0.465 ;
        RECT  7.225 -0.235 7.675 0.235 ;
        RECT  6.815 -0.235 7.225 0.465 ;
        RECT  3.945 -0.235 6.815 0.235 ;
        RECT  3.605 -0.235 3.945 0.465 ;
        RECT  1.265 -0.235 3.605 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.805 3.685 19.040 4.155 ;
        RECT  18.575 2.255 18.805 4.155 ;
        RECT  17.420 3.685 18.575 4.155 ;
        RECT  17.080 3.250 17.420 4.155 ;
        RECT  15.860 3.685 17.080 4.155 ;
        RECT  15.520 3.455 15.860 4.155 ;
        RECT  14.345 3.685 15.520 4.155 ;
        RECT  14.005 3.455 14.345 4.155 ;
        RECT  11.650 3.685 14.005 4.155 ;
        RECT  11.290 3.190 11.650 4.155 ;
        RECT  8.230 3.685 11.290 4.155 ;
        RECT  7.890 3.455 8.230 4.155 ;
        RECT  7.170 3.685 7.890 4.155 ;
        RECT  6.830 3.455 7.170 4.155 ;
        RECT  4.775 3.685 6.830 4.155 ;
        RECT  4.435 3.455 4.775 4.155 ;
        RECT  1.265 3.685 4.435 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.375 1.600 17.605 3.020 ;
        RECT  16.070 2.790 17.375 3.020 ;
        RECT  15.160 1.615 16.130 1.955 ;
        RECT  15.840 2.790 16.070 3.215 ;
        RECT  14.220 2.985 15.840 3.215 ;
        RECT  14.930 0.465 15.160 2.755 ;
        RECT  14.010 0.940 14.930 1.170 ;
        RECT  14.810 2.520 14.930 2.755 ;
        RECT  14.450 1.565 14.680 2.290 ;
        RECT  14.220 2.060 14.450 2.290 ;
        RECT  13.990 2.060 14.220 3.215 ;
        RECT  13.780 0.940 14.010 1.830 ;
        RECT  13.065 2.060 13.990 2.290 ;
        RECT  12.355 3.225 13.500 3.455 ;
        RECT  12.835 0.910 13.065 2.850 ;
        RECT  12.375 0.960 12.605 2.500 ;
        RECT  11.325 0.960 12.375 1.190 ;
        RECT  12.060 2.270 12.375 2.500 ;
        RECT  12.125 2.730 12.355 3.455 ;
        RECT  10.950 2.730 12.125 2.960 ;
        RECT  11.830 1.560 12.105 1.900 ;
        RECT  11.600 1.560 11.830 2.415 ;
        RECT  10.395 2.185 11.600 2.415 ;
        RECT  11.095 0.960 11.325 1.890 ;
        RECT  10.720 2.730 10.950 3.375 ;
        RECT  9.175 3.145 10.720 3.375 ;
        RECT  10.355 0.935 10.395 2.415 ;
        RECT  10.125 0.935 10.355 2.905 ;
        RECT  9.730 1.005 9.875 2.840 ;
        RECT  9.645 0.520 9.730 2.840 ;
        RECT  9.390 0.520 9.645 1.220 ;
        RECT  9.405 2.420 9.645 2.840 ;
        RECT  8.465 0.520 9.390 0.750 ;
        RECT  9.175 1.615 9.350 1.955 ;
        RECT  9.150 1.615 9.175 3.375 ;
        RECT  8.945 0.980 9.150 3.375 ;
        RECT  8.920 0.980 8.945 2.760 ;
        RECT  8.690 0.980 8.920 1.210 ;
        RECT  8.645 2.530 8.920 2.760 ;
        RECT  8.465 2.995 8.695 3.455 ;
        RECT  8.240 0.520 8.465 0.925 ;
        RECT  7.675 2.995 8.465 3.225 ;
        RECT  6.355 0.695 8.240 0.925 ;
        RECT  7.445 2.560 7.675 3.225 ;
        RECT  7.425 1.155 7.670 1.385 ;
        RECT  7.425 2.560 7.445 2.790 ;
        RECT  7.195 1.155 7.425 2.790 ;
        RECT  6.645 1.620 6.875 3.225 ;
        RECT  2.615 2.995 6.645 3.225 ;
        RECT  6.115 0.495 6.355 2.765 ;
        RECT  4.870 0.480 5.710 0.710 ;
        RECT  4.870 2.450 5.680 2.680 ;
        RECT  4.640 0.480 4.870 2.680 ;
        RECT  4.185 1.665 4.640 1.895 ;
        RECT  3.930 1.020 4.390 1.250 ;
        RECT  3.700 0.750 3.930 2.680 ;
        RECT  3.075 0.750 3.700 0.980 ;
        RECT  2.940 2.450 3.700 2.680 ;
        RECT  2.845 0.510 3.075 0.980 ;
        RECT  2.385 0.850 2.615 3.225 ;
        RECT  2.050 0.850 2.385 1.080 ;
        RECT  2.130 2.440 2.385 2.680 ;
        RECT  1.925 1.310 2.155 2.080 ;
        RECT  0.465 1.310 1.925 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKSND2BWP7T

MACRO SDFKSNQD0BWP7T
    CLASS CORE ;
    FOREIGN SDFKSNQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.210 5.460 2.150 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.560 16.660 2.975 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.680 3.420 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.760 8.260 2.710 ;
        RECT  7.740 1.760 7.980 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.845 -0.235 16.800 0.235 ;
        RECT  15.615 -0.235 15.845 0.910 ;
        RECT  14.420 -0.235 15.615 0.235 ;
        RECT  14.080 -0.235 14.420 0.720 ;
        RECT  11.640 -0.235 14.080 0.235 ;
        RECT  11.300 -0.235 11.640 0.730 ;
        RECT  8.015 -0.235 11.300 0.235 ;
        RECT  7.675 -0.235 8.015 0.465 ;
        RECT  7.225 -0.235 7.675 0.235 ;
        RECT  6.815 -0.235 7.225 0.465 ;
        RECT  3.945 -0.235 6.815 0.235 ;
        RECT  3.605 -0.235 3.945 0.465 ;
        RECT  1.265 -0.235 3.605 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.845 3.685 16.800 4.155 ;
        RECT  15.615 2.645 15.845 4.155 ;
        RECT  14.440 3.685 15.615 4.155 ;
        RECT  14.100 2.665 14.440 4.155 ;
        RECT  11.650 3.685 14.100 4.155 ;
        RECT  11.290 3.190 11.650 4.155 ;
        RECT  8.230 3.685 11.290 4.155 ;
        RECT  7.890 3.455 8.230 4.155 ;
        RECT  7.170 3.685 7.890 4.155 ;
        RECT  6.830 3.455 7.170 4.155 ;
        RECT  4.775 3.685 6.830 4.155 ;
        RECT  4.435 3.455 4.775 4.155 ;
        RECT  1.265 3.685 4.435 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.155 0.950 15.385 2.915 ;
        RECT  14.010 0.950 15.155 1.180 ;
        RECT  14.860 2.680 15.155 2.915 ;
        RECT  14.675 1.605 14.905 2.290 ;
        RECT  13.065 2.060 14.675 2.290 ;
        RECT  13.780 0.950 14.010 1.830 ;
        RECT  12.355 3.225 13.480 3.455 ;
        RECT  12.835 0.910 13.065 2.850 ;
        RECT  12.375 0.960 12.605 2.500 ;
        RECT  11.325 0.960 12.375 1.190 ;
        RECT  12.060 2.270 12.375 2.500 ;
        RECT  12.125 2.730 12.355 3.455 ;
        RECT  10.950 2.730 12.125 2.960 ;
        RECT  11.830 1.560 12.105 1.900 ;
        RECT  11.600 1.560 11.830 2.415 ;
        RECT  10.395 2.185 11.600 2.415 ;
        RECT  11.095 0.960 11.325 1.890 ;
        RECT  10.720 2.730 10.950 3.375 ;
        RECT  9.175 3.145 10.720 3.375 ;
        RECT  10.355 0.935 10.395 2.415 ;
        RECT  10.125 0.935 10.355 2.905 ;
        RECT  9.730 1.005 9.875 2.840 ;
        RECT  9.645 0.520 9.730 2.840 ;
        RECT  9.390 0.520 9.645 1.220 ;
        RECT  9.405 2.420 9.645 2.840 ;
        RECT  8.465 0.520 9.390 0.750 ;
        RECT  9.175 1.615 9.350 1.955 ;
        RECT  9.150 1.615 9.175 3.375 ;
        RECT  8.945 0.980 9.150 3.375 ;
        RECT  8.920 0.980 8.945 2.760 ;
        RECT  8.690 0.980 8.920 1.210 ;
        RECT  8.645 2.530 8.920 2.760 ;
        RECT  8.465 2.995 8.695 3.455 ;
        RECT  8.240 0.520 8.465 0.925 ;
        RECT  7.675 2.995 8.465 3.225 ;
        RECT  6.355 0.695 8.240 0.925 ;
        RECT  7.445 2.560 7.675 3.225 ;
        RECT  7.425 1.155 7.670 1.385 ;
        RECT  7.425 2.560 7.445 2.790 ;
        RECT  7.195 1.155 7.425 2.790 ;
        RECT  6.645 1.620 6.875 3.225 ;
        RECT  2.615 2.995 6.645 3.225 ;
        RECT  6.115 0.495 6.355 2.765 ;
        RECT  4.870 0.480 5.710 0.710 ;
        RECT  4.870 2.450 5.680 2.680 ;
        RECT  4.640 0.480 4.870 2.680 ;
        RECT  4.185 1.665 4.640 1.895 ;
        RECT  3.930 1.020 4.390 1.250 ;
        RECT  3.700 0.750 3.930 2.680 ;
        RECT  3.075 0.750 3.700 0.980 ;
        RECT  2.940 2.450 3.700 2.680 ;
        RECT  2.845 0.510 3.075 0.980 ;
        RECT  2.385 0.850 2.615 3.225 ;
        RECT  2.050 0.850 2.385 1.080 ;
        RECT  2.130 2.440 2.385 2.680 ;
        RECT  1.925 1.310 2.155 2.080 ;
        RECT  0.465 1.310 1.925 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKSNQD0BWP7T

MACRO SDFKSNQD1BWP7T
    CLASS CORE ;
    FOREIGN SDFKSNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.210 5.460 2.150 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.470 16.660 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.680 3.420 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.760 8.260 2.710 ;
        RECT  7.740 1.760 7.980 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.845 -0.235 16.800 0.235 ;
        RECT  15.615 -0.235 15.845 1.245 ;
        RECT  14.420 -0.235 15.615 0.235 ;
        RECT  14.080 -0.235 14.420 0.720 ;
        RECT  11.640 -0.235 14.080 0.235 ;
        RECT  11.300 -0.235 11.640 0.730 ;
        RECT  8.015 -0.235 11.300 0.235 ;
        RECT  7.675 -0.235 8.015 0.465 ;
        RECT  7.225 -0.235 7.675 0.235 ;
        RECT  6.815 -0.235 7.225 0.465 ;
        RECT  3.945 -0.235 6.815 0.235 ;
        RECT  3.605 -0.235 3.945 0.465 ;
        RECT  1.265 -0.235 3.605 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.845 3.685 16.800 4.155 ;
        RECT  15.615 2.255 15.845 4.155 ;
        RECT  14.440 3.685 15.615 4.155 ;
        RECT  14.100 2.665 14.440 4.155 ;
        RECT  11.650 3.685 14.100 4.155 ;
        RECT  11.290 3.190 11.650 4.155 ;
        RECT  8.230 3.685 11.290 4.155 ;
        RECT  7.890 3.455 8.230 4.155 ;
        RECT  7.170 3.685 7.890 4.155 ;
        RECT  6.830 3.455 7.170 4.155 ;
        RECT  4.775 3.685 6.830 4.155 ;
        RECT  4.435 3.455 4.775 4.155 ;
        RECT  1.265 3.685 4.435 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.155 0.950 15.385 2.915 ;
        RECT  14.010 0.950 15.155 1.180 ;
        RECT  14.860 2.680 15.155 2.915 ;
        RECT  14.675 1.605 14.905 2.290 ;
        RECT  13.065 2.060 14.675 2.290 ;
        RECT  13.780 0.950 14.010 1.830 ;
        RECT  12.355 3.225 13.480 3.455 ;
        RECT  12.835 0.910 13.065 2.850 ;
        RECT  12.375 0.960 12.605 2.500 ;
        RECT  11.325 0.960 12.375 1.190 ;
        RECT  12.060 2.270 12.375 2.500 ;
        RECT  12.125 2.730 12.355 3.455 ;
        RECT  10.950 2.730 12.125 2.960 ;
        RECT  11.830 1.560 12.105 1.900 ;
        RECT  11.600 1.560 11.830 2.415 ;
        RECT  10.395 2.185 11.600 2.415 ;
        RECT  11.095 0.960 11.325 1.890 ;
        RECT  10.720 2.730 10.950 3.375 ;
        RECT  9.175 3.145 10.720 3.375 ;
        RECT  10.355 0.935 10.395 2.415 ;
        RECT  10.125 0.935 10.355 2.905 ;
        RECT  9.730 1.000 9.875 2.840 ;
        RECT  9.645 0.520 9.730 2.840 ;
        RECT  9.390 0.520 9.645 1.220 ;
        RECT  9.405 2.420 9.645 2.840 ;
        RECT  8.465 0.520 9.390 0.750 ;
        RECT  9.175 1.615 9.350 1.955 ;
        RECT  9.150 1.615 9.175 3.375 ;
        RECT  8.945 0.980 9.150 3.375 ;
        RECT  8.920 0.980 8.945 2.760 ;
        RECT  8.690 0.980 8.920 1.210 ;
        RECT  8.645 2.530 8.920 2.760 ;
        RECT  8.465 2.995 8.695 3.455 ;
        RECT  8.240 0.520 8.465 0.925 ;
        RECT  7.675 2.995 8.465 3.225 ;
        RECT  6.355 0.695 8.240 0.925 ;
        RECT  7.445 2.560 7.675 3.225 ;
        RECT  7.425 1.155 7.670 1.385 ;
        RECT  7.425 2.560 7.445 2.790 ;
        RECT  7.195 1.155 7.425 2.790 ;
        RECT  6.645 1.620 6.875 3.225 ;
        RECT  2.615 2.995 6.645 3.225 ;
        RECT  6.115 0.495 6.355 2.765 ;
        RECT  4.870 0.480 5.710 0.710 ;
        RECT  4.870 2.450 5.680 2.680 ;
        RECT  4.640 0.480 4.870 2.680 ;
        RECT  4.185 1.665 4.640 1.895 ;
        RECT  3.930 1.020 4.390 1.250 ;
        RECT  3.700 0.750 3.930 2.680 ;
        RECT  3.075 0.750 3.700 0.980 ;
        RECT  2.940 2.450 3.700 2.680 ;
        RECT  2.845 0.510 3.075 0.980 ;
        RECT  2.385 0.850 2.615 3.225 ;
        RECT  2.050 0.850 2.385 1.080 ;
        RECT  2.130 2.440 2.385 2.680 ;
        RECT  1.925 1.310 2.155 2.080 ;
        RECT  0.465 1.310 1.925 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKSNQD1BWP7T

MACRO SDFKSNQD2BWP7T
    CLASS CORE ;
    FOREIGN SDFKSNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.360 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.125 1.210 5.460 2.150 ;
        END
    END SN
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.770 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4959 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.585 1.770 0.700 2.140 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.405 1.060 16.660 2.725 ;
        RECT  16.380 0.470 16.405 3.310 ;
        RECT  16.175 0.470 16.380 1.290 ;
        RECT  16.175 2.495 16.380 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.680 3.420 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.760 8.260 2.710 ;
        RECT  7.740 1.760 7.980 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.125 -0.235 17.360 0.235 ;
        RECT  16.895 -0.235 17.125 1.245 ;
        RECT  15.685 -0.235 16.895 0.235 ;
        RECT  15.455 -0.235 15.685 1.245 ;
        RECT  14.245 -0.235 15.455 0.235 ;
        RECT  13.905 -0.235 14.245 0.465 ;
        RECT  11.640 -0.235 13.905 0.235 ;
        RECT  11.300 -0.235 11.640 0.730 ;
        RECT  8.015 -0.235 11.300 0.235 ;
        RECT  7.675 -0.235 8.015 0.465 ;
        RECT  7.225 -0.235 7.675 0.235 ;
        RECT  6.815 -0.235 7.225 0.465 ;
        RECT  3.945 -0.235 6.815 0.235 ;
        RECT  3.605 -0.235 3.945 0.465 ;
        RECT  1.265 -0.235 3.605 0.235 ;
        RECT  0.885 -0.235 1.265 1.080 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.125 3.685 17.360 4.155 ;
        RECT  16.895 2.255 17.125 4.155 ;
        RECT  15.685 3.685 16.895 4.155 ;
        RECT  15.455 2.255 15.685 4.155 ;
        RECT  14.255 3.685 15.455 4.155 ;
        RECT  13.915 3.350 14.255 4.155 ;
        RECT  11.650 3.685 13.915 4.155 ;
        RECT  11.290 3.190 11.650 4.155 ;
        RECT  8.230 3.685 11.290 4.155 ;
        RECT  7.890 3.455 8.230 4.155 ;
        RECT  7.170 3.685 7.890 4.155 ;
        RECT  6.830 3.455 7.170 4.155 ;
        RECT  4.775 3.685 6.830 4.155 ;
        RECT  4.435 3.455 4.775 4.155 ;
        RECT  1.265 3.685 4.435 4.155 ;
        RECT  0.885 2.990 1.265 4.155 ;
        RECT  0.000 3.685 0.885 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.995 0.950 15.225 2.915 ;
        RECT  14.010 0.950 14.995 1.180 ;
        RECT  14.700 2.680 14.995 2.915 ;
        RECT  14.515 1.610 14.745 2.410 ;
        RECT  13.065 2.180 14.515 2.410 ;
        RECT  13.780 0.950 14.010 1.905 ;
        RECT  12.355 3.225 13.480 3.455 ;
        RECT  12.835 0.910 13.065 2.850 ;
        RECT  12.375 0.960 12.605 2.500 ;
        RECT  11.325 0.960 12.375 1.190 ;
        RECT  12.060 2.270 12.375 2.500 ;
        RECT  12.125 2.730 12.355 3.455 ;
        RECT  10.950 2.730 12.125 2.960 ;
        RECT  11.830 1.560 12.105 1.900 ;
        RECT  11.600 1.560 11.830 2.415 ;
        RECT  10.395 2.185 11.600 2.415 ;
        RECT  11.095 0.960 11.325 1.890 ;
        RECT  10.720 2.730 10.950 3.375 ;
        RECT  9.175 3.145 10.720 3.375 ;
        RECT  10.355 0.935 10.395 2.415 ;
        RECT  10.125 0.935 10.355 2.905 ;
        RECT  9.730 1.005 9.850 2.840 ;
        RECT  9.620 0.520 9.730 2.840 ;
        RECT  9.390 0.520 9.620 1.220 ;
        RECT  9.405 2.420 9.620 2.840 ;
        RECT  8.465 0.520 9.390 0.750 ;
        RECT  9.175 1.615 9.350 1.955 ;
        RECT  9.150 1.615 9.175 3.375 ;
        RECT  8.945 0.980 9.150 3.375 ;
        RECT  8.920 0.980 8.945 2.760 ;
        RECT  8.690 0.980 8.920 1.210 ;
        RECT  8.645 2.530 8.920 2.760 ;
        RECT  8.465 2.995 8.695 3.455 ;
        RECT  8.240 0.520 8.465 0.925 ;
        RECT  7.675 2.995 8.465 3.225 ;
        RECT  6.355 0.695 8.240 0.925 ;
        RECT  7.445 2.560 7.675 3.225 ;
        RECT  7.425 1.155 7.670 1.385 ;
        RECT  7.425 2.560 7.445 2.790 ;
        RECT  7.195 1.155 7.425 2.790 ;
        RECT  6.645 1.620 6.875 3.225 ;
        RECT  2.615 2.995 6.645 3.225 ;
        RECT  6.115 0.495 6.355 2.765 ;
        RECT  4.870 0.480 5.710 0.710 ;
        RECT  4.870 2.450 5.680 2.680 ;
        RECT  4.640 0.480 4.870 2.680 ;
        RECT  4.185 1.665 4.640 1.895 ;
        RECT  3.930 1.020 4.390 1.250 ;
        RECT  3.700 0.750 3.930 2.680 ;
        RECT  3.075 0.750 3.700 0.980 ;
        RECT  2.940 2.450 3.700 2.680 ;
        RECT  2.845 0.510 3.075 0.980 ;
        RECT  2.385 0.850 2.615 3.225 ;
        RECT  2.050 0.850 2.385 1.080 ;
        RECT  2.130 2.440 2.385 2.680 ;
        RECT  1.925 1.310 2.155 2.080 ;
        RECT  0.465 1.310 1.925 1.540 ;
        RECT  0.350 2.980 0.520 3.220 ;
        RECT  0.350 0.780 0.465 1.540 ;
        RECT  0.235 0.780 0.350 3.220 ;
        RECT  0.120 1.310 0.235 3.220 ;
    END
END SDFKSNQD2BWP7T

MACRO SDFNCND0BWP7T
    CLASS CORE ;
    FOREIGN SDFNCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.150 15.540 2.560 ;
        RECT  15.125 1.150 15.260 1.380 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.585 15.125 1.380 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.590 16.660 2.705 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.600 3.475 1.940 ;
        RECT  2.940 1.600 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.370 1.615 4.620 1.955 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.225 11.925 3.455 ;
        RECT  10.805 2.730 11.035 3.455 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.885 ;
        RECT  12.255 -0.235 15.560 0.235 ;
        RECT  11.915 -0.235 12.255 0.465 ;
        RECT  9.085 -0.235 11.915 0.235 ;
        RECT  8.745 -0.235 9.085 1.100 ;
        RECT  4.045 -0.235 8.745 0.235 ;
        RECT  3.705 -0.235 4.045 0.465 ;
        RECT  1.240 -0.235 3.705 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.820 3.685 16.800 4.155 ;
        RECT  15.480 3.455 15.820 4.155 ;
        RECT  14.640 3.685 15.480 4.155 ;
        RECT  14.300 3.455 14.640 4.155 ;
        RECT  13.110 3.685 14.300 4.155 ;
        RECT  12.770 3.190 13.110 4.155 ;
        RECT  10.575 3.685 12.770 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.875 3.685 10.235 4.155 ;
        RECT  4.535 3.455 4.875 4.155 ;
        RECT  3.840 3.685 4.535 4.155 ;
        RECT  3.500 3.455 3.840 4.155 ;
        RECT  1.240 3.685 3.500 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  14.575 2.790 15.855 3.020 ;
        RECT  12.850 0.465 14.660 0.695 ;
        RECT  14.345 0.990 14.575 3.020 ;
        RECT  13.455 0.990 14.345 1.220 ;
        RECT  13.820 2.490 14.345 2.720 ;
        RECT  13.835 1.565 14.065 2.260 ;
        RECT  13.015 2.030 13.835 2.260 ;
        RECT  13.590 2.490 13.820 3.335 ;
        RECT  13.225 0.990 13.455 1.760 ;
        RECT  12.280 1.530 13.225 1.760 ;
        RECT  12.785 2.030 13.015 2.960 ;
        RECT  12.620 0.465 12.850 1.220 ;
        RECT  11.495 2.730 12.785 2.960 ;
        RECT  12.000 0.990 12.620 1.220 ;
        RECT  12.000 2.270 12.270 2.500 ;
        RECT  11.770 0.990 12.000 2.500 ;
        RECT  11.015 0.990 11.770 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.785 1.330 9.810 1.560 ;
        RECT  9.555 0.870 9.785 1.560 ;
        RECT  8.805 1.330 9.555 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.300 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  5.360 0.465 7.715 0.695 ;
        RECT  7.100 0.935 7.300 2.230 ;
        RECT  7.070 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.070 3.085 ;
        RECT  6.380 0.925 6.605 2.505 ;
        RECT  6.375 0.925 6.380 3.225 ;
        RECT  6.255 0.925 6.375 1.155 ;
        RECT  6.150 2.275 6.375 3.225 ;
        RECT  2.600 2.995 6.150 3.225 ;
        RECT  5.840 1.615 6.100 1.955 ;
        RECT  5.610 0.925 5.840 2.765 ;
        RECT  5.290 2.535 5.610 2.765 ;
        RECT  5.130 0.465 5.360 1.970 ;
        RECT  4.030 0.975 5.130 1.205 ;
        RECT  4.030 2.425 4.260 2.765 ;
        RECT  3.800 0.975 4.030 2.765 ;
        RECT  2.480 1.075 2.600 3.225 ;
        RECT  2.370 0.465 2.480 3.225 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFNCND0BWP7T

MACRO SDFNCND1BWP7T
    CLASS CORE ;
    FOREIGN SDFNCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.9672 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.075 15.540 2.560 ;
        RECT  15.125 1.075 15.260 1.305 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.480 15.125 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.470 16.660 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.600 3.475 1.940 ;
        RECT  2.940 1.600 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.370 1.615 4.620 1.955 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.225 11.925 3.455 ;
        RECT  10.805 2.730 11.035 3.455 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.810 ;
        RECT  12.255 -0.235 15.560 0.235 ;
        RECT  11.915 -0.235 12.255 0.465 ;
        RECT  9.085 -0.235 11.915 0.235 ;
        RECT  8.745 -0.235 9.085 1.100 ;
        RECT  4.045 -0.235 8.745 0.235 ;
        RECT  3.705 -0.235 4.045 0.465 ;
        RECT  1.240 -0.235 3.705 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 3.685 16.800 4.155 ;
        RECT  15.560 3.250 15.900 4.155 ;
        RECT  14.640 3.685 15.560 4.155 ;
        RECT  14.300 3.455 14.640 4.155 ;
        RECT  13.110 3.685 14.300 4.155 ;
        RECT  12.770 3.190 13.110 4.155 ;
        RECT  10.575 3.685 12.770 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.875 3.685 10.235 4.155 ;
        RECT  4.535 3.455 4.875 4.155 ;
        RECT  3.840 3.685 4.535 4.155 ;
        RECT  3.500 3.455 3.840 4.155 ;
        RECT  1.240 3.685 3.500 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  14.575 2.790 15.855 3.020 ;
        RECT  12.850 0.465 14.660 0.695 ;
        RECT  14.345 1.020 14.575 3.020 ;
        RECT  13.455 1.020 14.345 1.250 ;
        RECT  13.820 2.565 14.345 2.795 ;
        RECT  13.835 1.565 14.065 2.260 ;
        RECT  13.015 2.030 13.835 2.260 ;
        RECT  13.590 2.565 13.820 3.375 ;
        RECT  13.225 1.020 13.455 1.760 ;
        RECT  12.280 1.530 13.225 1.760 ;
        RECT  12.785 2.030 13.015 2.960 ;
        RECT  12.620 0.465 12.850 1.220 ;
        RECT  11.495 2.730 12.785 2.960 ;
        RECT  12.000 0.990 12.620 1.220 ;
        RECT  12.000 2.270 12.270 2.500 ;
        RECT  11.770 0.990 12.000 2.500 ;
        RECT  11.015 0.990 11.770 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.785 1.330 9.810 1.560 ;
        RECT  9.555 0.870 9.785 1.560 ;
        RECT  8.805 1.330 9.555 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.300 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  5.360 0.465 7.715 0.695 ;
        RECT  7.100 0.935 7.300 2.230 ;
        RECT  7.070 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.070 3.085 ;
        RECT  6.380 0.925 6.605 2.505 ;
        RECT  6.375 0.925 6.380 3.225 ;
        RECT  6.255 0.925 6.375 1.155 ;
        RECT  6.150 2.275 6.375 3.225 ;
        RECT  2.600 2.995 6.150 3.225 ;
        RECT  5.840 1.615 6.100 1.955 ;
        RECT  5.610 0.925 5.840 2.765 ;
        RECT  5.290 2.535 5.610 2.765 ;
        RECT  5.130 0.465 5.360 1.970 ;
        RECT  4.030 0.975 5.130 1.205 ;
        RECT  4.030 2.425 4.260 2.765 ;
        RECT  3.800 0.975 4.030 2.765 ;
        RECT  2.480 1.075 2.600 3.225 ;
        RECT  2.370 0.465 2.480 3.225 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFNCND1BWP7T

MACRO SDFNCND2BWP7T
    CLASS CORE ;
    FOREIGN SDFNCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.240 0.465 15.585 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 1.055 17.220 2.690 ;
        RECT  16.940 0.465 16.965 3.310 ;
        RECT  16.730 0.465 16.940 1.285 ;
        RECT  16.735 2.460 16.940 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.600 3.475 1.940 ;
        RECT  2.940 1.600 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.615 4.900 2.710 ;
        RECT  4.370 1.615 4.620 1.955 ;
        END
    END CPN
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.035 3.190 11.765 3.420 ;
        RECT  10.805 2.730 11.035 3.420 ;
        RECT  9.870 2.730 10.805 2.960 ;
        RECT  9.640 2.730 9.870 3.270 ;
        RECT  7.895 2.940 9.640 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 -0.235 17.920 0.235 ;
        RECT  17.455 -0.235 17.685 1.245 ;
        RECT  16.300 -0.235 17.455 0.235 ;
        RECT  15.960 -0.235 16.300 1.180 ;
        RECT  14.820 -0.235 15.960 0.235 ;
        RECT  14.480 -0.235 14.820 0.465 ;
        RECT  12.890 -0.235 14.480 0.235 ;
        RECT  12.550 -0.235 12.890 0.465 ;
        RECT  9.085 -0.235 12.550 0.235 ;
        RECT  8.745 -0.235 9.085 1.100 ;
        RECT  4.045 -0.235 8.745 0.235 ;
        RECT  3.705 -0.235 4.045 0.465 ;
        RECT  1.240 -0.235 3.705 0.235 ;
        RECT  0.900 -0.235 1.240 0.880 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 3.685 17.920 4.155 ;
        RECT  17.455 2.255 17.685 4.155 ;
        RECT  16.300 3.685 17.455 4.155 ;
        RECT  15.960 3.250 16.300 4.155 ;
        RECT  14.705 3.685 15.960 4.155 ;
        RECT  14.365 3.250 14.705 4.155 ;
        RECT  13.105 3.685 14.365 4.155 ;
        RECT  12.765 3.190 13.105 4.155 ;
        RECT  10.575 3.685 12.765 4.155 ;
        RECT  10.235 3.190 10.575 4.155 ;
        RECT  4.875 3.685 10.235 4.155 ;
        RECT  4.535 3.455 4.875 4.155 ;
        RECT  3.840 3.685 4.535 4.155 ;
        RECT  3.500 3.455 3.840 4.155 ;
        RECT  1.240 3.685 3.500 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.255 1.600 16.485 3.020 ;
        RECT  14.480 2.790 16.255 3.020 ;
        RECT  14.770 0.695 15.000 1.940 ;
        RECT  12.075 0.695 14.770 0.925 ;
        RECT  14.250 1.155 14.480 3.020 ;
        RECT  13.035 1.155 14.250 1.385 ;
        RECT  13.825 2.540 14.250 2.770 ;
        RECT  13.720 1.670 13.950 2.260 ;
        RECT  13.595 2.540 13.825 3.370 ;
        RECT  13.055 2.030 13.720 2.260 ;
        RECT  12.825 2.030 13.055 2.960 ;
        RECT  12.805 1.155 13.035 1.750 ;
        RECT  11.495 2.730 12.825 2.960 ;
        RECT  12.305 1.520 12.805 1.750 ;
        RECT  12.075 2.270 12.270 2.500 ;
        RECT  11.845 0.465 12.075 2.500 ;
        RECT  10.970 0.990 11.845 1.220 ;
        RECT  11.265 1.615 11.495 2.960 ;
        RECT  10.720 1.615 11.265 1.845 ;
        RECT  10.490 0.985 10.720 1.845 ;
        RECT  10.040 2.270 10.640 2.500 ;
        RECT  10.250 0.985 10.490 1.220 ;
        RECT  9.810 1.330 10.040 2.500 ;
        RECT  9.785 1.330 9.810 1.560 ;
        RECT  9.555 0.870 9.785 1.560 ;
        RECT  8.805 1.330 9.555 1.560 ;
        RECT  9.165 1.790 9.505 2.230 ;
        RECT  7.655 2.460 9.315 2.690 ;
        RECT  7.300 2.000 9.165 2.230 ;
        RECT  8.465 1.330 8.805 1.770 ;
        RECT  5.360 0.465 7.715 0.695 ;
        RECT  7.100 0.935 7.300 2.230 ;
        RECT  7.070 0.935 7.100 3.085 ;
        RECT  6.865 2.000 7.070 3.085 ;
        RECT  6.380 0.925 6.605 2.505 ;
        RECT  6.375 0.925 6.380 3.225 ;
        RECT  6.255 0.925 6.375 1.155 ;
        RECT  6.150 2.275 6.375 3.225 ;
        RECT  2.600 2.995 6.150 3.225 ;
        RECT  5.840 1.615 6.100 1.955 ;
        RECT  5.610 0.925 5.840 2.765 ;
        RECT  5.290 2.535 5.610 2.765 ;
        RECT  5.130 0.465 5.360 1.970 ;
        RECT  4.030 0.975 5.130 1.205 ;
        RECT  4.030 2.425 4.260 2.765 ;
        RECT  3.800 0.975 4.030 2.765 ;
        RECT  2.480 1.075 2.600 3.225 ;
        RECT  2.370 0.465 2.480 3.225 ;
        RECT  2.250 0.465 2.370 1.280 ;
        RECT  2.090 2.770 2.370 3.000 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFNCND2BWP7T

MACRO SDFND0BWP7T
    CLASS CORE ;
    FOREIGN SDFND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.075 13.300 2.560 ;
        RECT  12.885 1.075 13.020 1.305 ;
        RECT  12.600 2.330 13.020 2.560 ;
        RECT  12.655 0.520 12.885 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.510 14.420 2.715 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.670 3.450 2.010 ;
        RECT  2.940 1.670 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.365 1.760 4.620 2.105 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.660 0.810 ;
        RECT  10.530 -0.235 13.320 0.235 ;
        RECT  10.190 -0.235 10.530 0.465 ;
        RECT  8.510 -0.235 10.190 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.795 -0.235 4.575 0.235 ;
        RECT  3.455 -0.235 3.795 0.465 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.730 3.685 14.560 4.155 ;
        RECT  13.390 3.365 13.730 4.155 ;
        RECT  11.430 3.685 13.390 4.155 ;
        RECT  11.090 3.385 11.430 4.155 ;
        RECT  8.520 3.685 11.090 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.860 3.685 8.160 4.155 ;
        RECT  4.520 3.455 4.860 4.155 ;
        RECT  3.790 3.685 4.520 4.155 ;
        RECT  3.450 3.455 3.790 4.155 ;
        RECT  1.240 3.685 3.450 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.020 ;
        RECT  12.370 2.790 13.615 3.020 ;
        RECT  10.990 0.465 12.420 0.695 ;
        RECT  12.140 1.020 12.370 3.020 ;
        RECT  11.450 1.020 12.140 1.250 ;
        RECT  11.900 2.540 12.140 2.775 ;
        RECT  11.680 1.565 11.910 2.310 ;
        RECT  11.450 2.080 11.680 2.310 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  11.220 2.080 11.450 2.995 ;
        RECT  10.735 1.600 11.220 1.830 ;
        RECT  9.935 2.765 11.220 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.500 2.300 10.770 2.530 ;
        RECT  10.500 0.990 10.760 1.220 ;
        RECT  10.270 0.990 10.500 2.530 ;
        RECT  9.225 3.225 10.480 3.455 ;
        RECT  9.705 0.910 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.455 ;
        RECT  5.320 3.225 7.520 3.455 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.380 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.640 6.085 1.980 ;
        RECT  5.615 0.925 5.845 2.720 ;
        RECT  5.275 2.490 5.615 2.720 ;
        RECT  5.150 0.465 5.380 0.925 ;
        RECT  5.130 1.155 5.360 2.090 ;
        RECT  5.090 2.960 5.320 3.455 ;
        RECT  2.655 0.695 5.150 0.925 ;
        RECT  3.990 1.155 5.130 1.385 ;
        RECT  4.300 2.960 5.090 3.190 ;
        RECT  4.070 2.560 4.300 3.190 ;
        RECT  3.990 2.560 4.070 2.790 ;
        RECT  3.760 1.155 3.990 2.790 ;
        RECT  2.460 0.695 2.655 2.780 ;
        RECT  2.425 0.695 2.460 3.355 ;
        RECT  2.195 0.695 2.425 0.925 ;
        RECT  2.230 2.545 2.425 3.355 ;
        RECT  2.025 1.780 2.190 2.010 ;
        RECT  1.795 1.130 2.025 2.010 ;
        RECT  0.465 1.130 1.795 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFND0BWP7T

MACRO SDFND1BWP7T
    CLASS CORE ;
    FOREIGN SDFND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.020 1.075 13.300 2.560 ;
        RECT  12.885 1.075 13.020 1.305 ;
        RECT  12.600 2.330 13.020 2.560 ;
        RECT  12.655 0.480 12.885 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.090 0.470 14.420 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.670 3.450 2.010 ;
        RECT  2.940 1.670 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.365 1.760 4.620 2.105 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 -0.235 14.560 0.235 ;
        RECT  13.320 -0.235 13.660 0.810 ;
        RECT  10.530 -0.235 13.320 0.235 ;
        RECT  10.190 -0.235 10.530 0.465 ;
        RECT  8.510 -0.235 10.190 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.795 -0.235 4.575 0.235 ;
        RECT  3.455 -0.235 3.795 0.465 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.660 3.685 14.560 4.155 ;
        RECT  13.320 3.250 13.660 4.155 ;
        RECT  11.520 3.685 13.320 4.155 ;
        RECT  11.180 3.250 11.520 4.155 ;
        RECT  8.520 3.685 11.180 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.860 3.685 8.160 4.155 ;
        RECT  4.520 3.455 4.860 4.155 ;
        RECT  3.790 3.685 4.520 4.155 ;
        RECT  3.450 3.455 3.790 4.155 ;
        RECT  1.240 3.685 3.450 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.600 13.845 3.020 ;
        RECT  12.370 2.790 13.615 3.020 ;
        RECT  10.990 0.465 12.420 0.695 ;
        RECT  12.185 1.020 12.370 3.020 ;
        RECT  12.140 1.020 12.185 3.380 ;
        RECT  11.450 1.020 12.140 1.250 ;
        RECT  11.955 2.565 12.140 3.380 ;
        RECT  11.680 1.565 11.910 2.310 ;
        RECT  11.450 2.080 11.680 2.310 ;
        RECT  11.220 1.020 11.450 1.830 ;
        RECT  11.220 2.080 11.450 2.995 ;
        RECT  10.735 1.600 11.220 1.830 ;
        RECT  9.935 2.765 11.220 2.995 ;
        RECT  10.760 0.465 10.990 1.220 ;
        RECT  10.500 2.300 10.770 2.530 ;
        RECT  10.500 0.990 10.760 1.220 ;
        RECT  10.270 0.990 10.500 2.530 ;
        RECT  9.225 3.225 10.480 3.455 ;
        RECT  9.705 0.910 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.455 ;
        RECT  5.320 3.225 7.520 3.455 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.380 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.640 6.085 1.980 ;
        RECT  5.615 0.925 5.845 2.720 ;
        RECT  5.275 2.490 5.615 2.720 ;
        RECT  5.150 0.465 5.380 0.925 ;
        RECT  5.130 1.155 5.360 2.090 ;
        RECT  5.090 2.960 5.320 3.455 ;
        RECT  2.655 0.695 5.150 0.925 ;
        RECT  3.990 1.155 5.130 1.385 ;
        RECT  4.300 2.960 5.090 3.190 ;
        RECT  4.070 2.560 4.300 3.190 ;
        RECT  3.990 2.560 4.070 2.790 ;
        RECT  3.760 1.155 3.990 2.790 ;
        RECT  2.460 0.695 2.655 2.780 ;
        RECT  2.425 0.695 2.460 3.355 ;
        RECT  2.195 0.695 2.425 0.925 ;
        RECT  2.230 2.545 2.425 3.355 ;
        RECT  2.025 1.780 2.190 2.010 ;
        RECT  1.795 1.130 2.025 2.010 ;
        RECT  0.465 1.130 1.795 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFND1BWP7T

MACRO SDFND2BWP7T
    CLASS CORE ;
    FOREIGN SDFND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.560 0.465 13.905 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.055 15.540 2.690 ;
        RECT  15.260 0.465 15.285 3.310 ;
        RECT  15.050 0.465 15.260 1.285 ;
        RECT  15.055 2.460 15.260 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.670 3.450 2.010 ;
        RECT  2.940 1.670 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.365 1.760 4.620 2.105 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.245 ;
        RECT  14.620 -0.235 15.775 0.235 ;
        RECT  14.280 -0.235 14.620 1.180 ;
        RECT  13.140 -0.235 14.280 0.235 ;
        RECT  12.800 -0.235 13.140 0.465 ;
        RECT  11.525 -0.235 12.800 0.235 ;
        RECT  11.185 -0.235 11.525 0.465 ;
        RECT  8.510 -0.235 11.185 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.795 -0.235 4.575 0.235 ;
        RECT  3.455 -0.235 3.795 0.465 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.255 16.005 4.155 ;
        RECT  14.620 3.685 15.775 4.155 ;
        RECT  14.280 3.250 14.620 4.155 ;
        RECT  13.105 3.685 14.280 4.155 ;
        RECT  12.765 3.250 13.105 4.155 ;
        RECT  11.575 3.685 12.765 4.155 ;
        RECT  11.235 3.250 11.575 4.155 ;
        RECT  8.520 3.685 11.235 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.860 3.685 8.160 4.155 ;
        RECT  4.520 3.455 4.860 4.155 ;
        RECT  3.790 3.685 4.520 4.155 ;
        RECT  3.450 3.455 3.790 4.155 ;
        RECT  1.240 3.685 3.450 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.575 1.600 14.805 3.010 ;
        RECT  12.555 2.780 14.575 3.010 ;
        RECT  13.090 0.695 13.320 1.940 ;
        RECT  10.990 0.695 13.090 0.925 ;
        RECT  12.325 1.155 12.555 3.010 ;
        RECT  11.505 1.155 12.325 1.385 ;
        RECT  12.285 2.565 12.325 3.010 ;
        RECT  12.055 2.565 12.285 3.380 ;
        RECT  11.800 1.675 12.030 2.310 ;
        RECT  11.530 2.080 11.800 2.310 ;
        RECT  11.300 2.080 11.530 2.995 ;
        RECT  11.275 1.155 11.505 1.830 ;
        RECT  9.935 2.765 11.300 2.995 ;
        RECT  10.725 1.600 11.275 1.830 ;
        RECT  10.760 0.695 10.990 1.220 ;
        RECT  10.460 2.300 10.770 2.530 ;
        RECT  10.460 0.990 10.760 1.220 ;
        RECT  10.230 0.990 10.460 2.530 ;
        RECT  9.225 3.225 10.425 3.455 ;
        RECT  9.705 0.910 9.935 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.455 ;
        RECT  5.320 3.225 7.520 3.455 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.380 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.640 6.085 1.980 ;
        RECT  5.615 0.925 5.845 2.720 ;
        RECT  5.275 2.490 5.615 2.720 ;
        RECT  5.150 0.465 5.380 0.925 ;
        RECT  5.130 1.155 5.360 2.090 ;
        RECT  5.090 2.960 5.320 3.455 ;
        RECT  2.655 0.695 5.150 0.925 ;
        RECT  3.990 1.155 5.130 1.385 ;
        RECT  4.300 2.960 5.090 3.190 ;
        RECT  4.070 2.560 4.300 3.190 ;
        RECT  3.990 2.560 4.070 2.790 ;
        RECT  3.760 1.155 3.990 2.790 ;
        RECT  2.460 0.695 2.655 2.780 ;
        RECT  2.425 0.695 2.460 3.355 ;
        RECT  2.195 0.695 2.425 0.925 ;
        RECT  2.230 2.545 2.425 3.355 ;
        RECT  2.025 1.780 2.190 2.010 ;
        RECT  1.795 1.130 2.025 2.010 ;
        RECT  0.465 1.130 1.795 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFND2BWP7T

MACRO SDFNSND0BWP7T
    CLASS CORE ;
    FOREIGN SDFNSND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.715 2.940 12.055 3.370 ;
        RECT  10.485 2.940 11.715 3.220 ;
        RECT  10.255 2.730 10.485 3.220 ;
        RECT  8.730 2.730 10.255 2.960 ;
        RECT  8.500 2.730 8.730 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.565 16.660 2.720 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.120 15.540 2.660 ;
        RECT  15.125 1.120 15.260 1.350 ;
        RECT  14.840 2.430 15.260 2.660 ;
        RECT  14.895 0.560 15.125 1.350 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.660 3.530 1.890 ;
        RECT  2.940 1.660 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 1.770 5.460 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.860 ;
        RECT  13.565 -0.235 15.560 0.235 ;
        RECT  13.225 -0.235 13.565 0.860 ;
        RECT  8.650 -0.235 13.225 0.235 ;
        RECT  8.310 -0.235 8.650 0.960 ;
        RECT  3.885 -0.235 8.310 0.235 ;
        RECT  3.545 -0.235 3.885 0.465 ;
        RECT  1.240 -0.235 3.545 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.830 3.685 16.800 4.155 ;
        RECT  15.490 3.455 15.830 4.155 ;
        RECT  13.715 3.685 15.490 4.155 ;
        RECT  13.375 3.455 13.715 4.155 ;
        RECT  12.690 3.685 13.375 4.155 ;
        RECT  12.350 3.450 12.690 4.155 ;
        RECT  9.920 3.685 12.350 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.875 3.685 7.980 4.155 ;
        RECT  4.535 3.455 4.875 4.155 ;
        RECT  3.825 3.685 4.535 4.155 ;
        RECT  3.485 3.455 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.410 16.085 3.225 ;
        RECT  13.325 2.995 15.855 3.225 ;
        RECT  14.610 1.635 15.030 1.865 ;
        RECT  14.425 0.630 14.610 2.230 ;
        RECT  14.380 0.630 14.425 2.765 ;
        RECT  13.990 0.630 14.380 0.860 ;
        RECT  14.195 2.000 14.380 2.765 ;
        RECT  13.080 2.000 14.195 2.230 ;
        RECT  13.805 1.205 14.035 1.750 ;
        RECT  12.800 1.205 13.805 1.435 ;
        RECT  13.090 2.465 13.325 3.225 ;
        RECT  11.845 2.465 13.090 2.695 ;
        RECT  12.740 1.780 13.080 2.230 ;
        RECT  12.570 0.465 12.800 1.435 ;
        RECT  10.580 0.465 12.570 0.695 ;
        RECT  11.845 0.990 12.170 1.220 ;
        RECT  11.615 0.990 11.845 2.695 ;
        RECT  11.015 0.990 11.615 1.220 ;
        RECT  10.895 1.615 11.125 2.585 ;
        RECT  10.580 1.615 10.895 1.845 ;
        RECT  10.350 0.465 10.580 1.845 ;
        RECT  10.120 2.270 10.460 2.500 ;
        RECT  9.890 0.935 10.120 2.500 ;
        RECT  9.510 0.935 9.890 1.165 ;
        RECT  8.195 2.270 9.890 2.500 ;
        RECT  8.965 1.640 9.610 1.870 ;
        RECT  8.735 1.190 8.965 1.870 ;
        RECT  7.220 1.190 8.735 1.420 ;
        RECT  7.965 1.650 8.195 2.500 ;
        RECT  4.735 0.465 7.700 0.695 ;
        RECT  7.100 0.990 7.220 1.420 ;
        RECT  6.870 0.990 7.100 3.085 ;
        RECT  6.380 0.925 6.600 2.505 ;
        RECT  6.370 0.925 6.380 3.225 ;
        RECT  6.150 0.925 6.370 1.155 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  2.600 2.995 6.150 3.225 ;
        RECT  5.920 1.605 6.100 1.945 ;
        RECT  5.690 1.005 5.920 2.765 ;
        RECT  5.290 1.005 5.690 1.235 ;
        RECT  5.290 2.535 5.690 2.765 ;
        RECT  4.505 0.465 4.735 1.210 ;
        RECT  4.065 0.980 4.505 1.210 ;
        RECT  4.065 2.535 4.315 2.765 ;
        RECT  3.835 0.980 4.065 2.765 ;
        RECT  2.480 1.085 2.600 3.225 ;
        RECT  2.370 0.465 2.480 3.225 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFNSND0BWP7T

MACRO SDFNSND1BWP7T
    CLASS CORE ;
    FOREIGN SDFNSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.715 2.940 12.055 3.370 ;
        RECT  10.485 2.940 11.715 3.220 ;
        RECT  10.255 2.730 10.485 3.220 ;
        RECT  8.730 2.730 10.255 2.960 ;
        RECT  8.500 2.730 8.730 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.470 16.660 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.075 15.540 2.560 ;
        RECT  15.125 1.075 15.260 1.305 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.465 15.125 1.305 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.660 3.530 1.890 ;
        RECT  2.940 1.660 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 1.770 5.460 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.810 ;
        RECT  13.565 -0.235 15.560 0.235 ;
        RECT  13.225 -0.235 13.565 0.930 ;
        RECT  8.650 -0.235 13.225 0.235 ;
        RECT  8.310 -0.235 8.650 0.960 ;
        RECT  3.885 -0.235 8.310 0.235 ;
        RECT  3.545 -0.235 3.885 0.465 ;
        RECT  1.240 -0.235 3.545 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 3.685 16.800 4.155 ;
        RECT  15.560 3.250 15.900 4.155 ;
        RECT  13.715 3.685 15.560 4.155 ;
        RECT  13.375 3.455 13.715 4.155 ;
        RECT  12.690 3.685 13.375 4.155 ;
        RECT  12.350 3.450 12.690 4.155 ;
        RECT  9.920 3.685 12.350 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.875 3.685 7.980 4.155 ;
        RECT  4.535 3.455 4.875 4.155 ;
        RECT  3.825 3.685 4.535 4.155 ;
        RECT  3.485 3.455 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  15.085 2.790 15.855 3.020 ;
        RECT  14.855 2.790 15.085 3.225 ;
        RECT  14.610 1.635 15.030 1.865 ;
        RECT  13.325 2.995 14.855 3.225 ;
        RECT  14.425 0.680 14.610 2.230 ;
        RECT  14.380 0.680 14.425 2.765 ;
        RECT  13.990 0.680 14.380 0.910 ;
        RECT  14.195 2.000 14.380 2.765 ;
        RECT  13.080 2.000 14.195 2.230 ;
        RECT  13.745 1.205 14.090 1.770 ;
        RECT  12.800 1.205 13.745 1.435 ;
        RECT  13.090 2.465 13.325 3.225 ;
        RECT  11.845 2.465 13.090 2.695 ;
        RECT  12.740 1.780 13.080 2.230 ;
        RECT  12.570 0.465 12.800 1.435 ;
        RECT  10.580 0.465 12.570 0.695 ;
        RECT  11.845 0.990 12.170 1.220 ;
        RECT  11.615 0.990 11.845 2.695 ;
        RECT  11.015 0.990 11.615 1.220 ;
        RECT  10.895 1.615 11.125 2.585 ;
        RECT  10.580 1.615 10.895 1.845 ;
        RECT  10.350 0.465 10.580 1.845 ;
        RECT  10.120 2.270 10.460 2.500 ;
        RECT  9.890 0.935 10.120 2.500 ;
        RECT  9.510 0.935 9.890 1.165 ;
        RECT  8.195 2.270 9.890 2.500 ;
        RECT  8.965 1.640 9.610 1.870 ;
        RECT  8.735 1.190 8.965 1.870 ;
        RECT  7.220 1.190 8.735 1.420 ;
        RECT  7.965 1.650 8.195 2.500 ;
        RECT  4.735 0.465 7.700 0.695 ;
        RECT  7.100 0.990 7.220 1.420 ;
        RECT  6.870 0.990 7.100 3.085 ;
        RECT  6.380 0.925 6.600 2.505 ;
        RECT  6.370 0.925 6.380 3.225 ;
        RECT  6.150 0.925 6.370 1.155 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  2.600 2.995 6.150 3.225 ;
        RECT  5.920 1.605 6.100 1.945 ;
        RECT  5.690 1.005 5.920 2.765 ;
        RECT  5.290 1.005 5.690 1.235 ;
        RECT  5.290 2.535 5.690 2.765 ;
        RECT  4.505 0.465 4.735 1.210 ;
        RECT  4.065 0.980 4.505 1.210 ;
        RECT  4.065 2.535 4.315 2.765 ;
        RECT  3.835 0.980 4.065 2.765 ;
        RECT  2.480 1.085 2.600 3.225 ;
        RECT  2.370 0.465 2.480 3.225 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFNSND1BWP7T

MACRO SDFNSND2BWP7T
    CLASS CORE ;
    FOREIGN SDFNSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.4491 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.205 3.225 13.620 3.455 ;
        RECT  11.975 2.935 12.205 3.455 ;
        RECT  10.380 2.935 11.975 3.220 ;
        RECT  10.150 2.730 10.380 3.220 ;
        RECT  8.730 2.730 10.150 2.960 ;
        RECT  8.500 2.730 8.730 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 1.055 17.220 2.690 ;
        RECT  16.940 0.465 16.965 3.310 ;
        RECT  16.730 0.465 16.940 1.285 ;
        RECT  16.735 2.460 16.940 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.240 0.545 15.585 2.530 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.660 3.530 1.890 ;
        RECT  2.940 1.660 3.220 2.710 ;
        END
    END D
    PIN CPN
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 1.770 5.460 2.150 ;
        END
    END CPN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 -0.235 17.920 0.235 ;
        RECT  17.455 -0.235 17.685 1.245 ;
        RECT  16.300 -0.235 17.455 0.235 ;
        RECT  15.960 -0.235 16.300 1.180 ;
        RECT  14.860 -0.235 15.960 0.235 ;
        RECT  14.520 -0.235 14.860 0.670 ;
        RECT  12.220 -0.235 14.520 0.235 ;
        RECT  11.990 -0.235 12.220 0.720 ;
        RECT  8.650 -0.235 11.990 0.235 ;
        RECT  8.310 -0.235 8.650 0.960 ;
        RECT  3.885 -0.235 8.310 0.235 ;
        RECT  3.545 -0.235 3.885 0.465 ;
        RECT  1.240 -0.235 3.545 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 3.685 17.920 4.155 ;
        RECT  17.455 2.255 17.685 4.155 ;
        RECT  16.300 3.685 17.455 4.155 ;
        RECT  15.960 3.250 16.300 4.155 ;
        RECT  14.860 3.685 15.960 4.155 ;
        RECT  14.520 3.250 14.860 4.155 ;
        RECT  11.745 3.685 14.520 4.155 ;
        RECT  11.405 3.450 11.745 4.155 ;
        RECT  9.920 3.685 11.405 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.875 3.685 7.980 4.155 ;
        RECT  4.535 3.455 4.875 4.155 ;
        RECT  3.825 3.685 4.535 4.155 ;
        RECT  3.485 3.455 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.255 1.600 16.485 2.990 ;
        RECT  15.010 2.760 16.255 2.990 ;
        RECT  14.780 0.900 15.010 2.990 ;
        RECT  13.870 0.900 14.780 1.130 ;
        RECT  12.665 2.760 14.780 2.990 ;
        RECT  13.285 1.620 14.550 1.960 ;
        RECT  13.640 0.465 13.870 1.130 ;
        RECT  13.355 0.465 13.640 0.695 ;
        RECT  13.055 0.945 13.285 2.530 ;
        RECT  12.655 0.945 13.055 1.175 ;
        RECT  12.910 2.300 13.055 2.530 ;
        RECT  12.285 1.540 12.800 1.770 ;
        RECT  12.435 2.300 12.665 2.990 ;
        RECT  11.585 2.300 12.435 2.530 ;
        RECT  12.055 0.950 12.285 1.770 ;
        RECT  11.750 0.950 12.055 1.180 ;
        RECT  11.520 0.465 11.750 1.180 ;
        RECT  11.355 1.410 11.585 2.530 ;
        RECT  10.530 0.465 11.520 0.695 ;
        RECT  11.290 1.410 11.355 1.640 ;
        RECT  11.060 0.935 11.290 1.640 ;
        RECT  10.880 2.245 11.125 2.585 ;
        RECT  10.650 1.810 10.880 2.585 ;
        RECT  10.530 1.810 10.650 2.040 ;
        RECT  10.300 0.465 10.530 2.040 ;
        RECT  10.070 2.270 10.420 2.500 ;
        RECT  9.840 0.935 10.070 2.500 ;
        RECT  9.495 0.935 9.840 1.165 ;
        RECT  8.195 2.270 9.840 2.500 ;
        RECT  8.965 1.640 9.610 1.870 ;
        RECT  8.735 1.190 8.965 1.870 ;
        RECT  7.220 1.190 8.735 1.420 ;
        RECT  7.965 1.650 8.195 2.500 ;
        RECT  4.735 0.465 7.700 0.695 ;
        RECT  7.100 0.990 7.220 1.420 ;
        RECT  6.870 0.990 7.100 3.085 ;
        RECT  6.380 0.925 6.600 2.505 ;
        RECT  6.370 0.925 6.380 3.225 ;
        RECT  6.150 0.925 6.370 1.155 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  2.600 2.995 6.150 3.225 ;
        RECT  5.920 1.605 6.100 1.945 ;
        RECT  5.690 1.005 5.920 2.765 ;
        RECT  5.290 1.005 5.690 1.235 ;
        RECT  5.290 2.535 5.690 2.765 ;
        RECT  4.505 0.465 4.735 1.210 ;
        RECT  4.065 0.980 4.505 1.210 ;
        RECT  4.065 2.535 4.315 2.765 ;
        RECT  3.835 0.980 4.065 2.765 ;
        RECT  2.480 1.085 2.600 3.225 ;
        RECT  2.370 0.465 2.480 3.225 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFNSND2BWP7T

MACRO SDFQD0BWP7T
    CLASS CORE ;
    FOREIGN SDFQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4824 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.970 0.585 13.300 3.195 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3474 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.680 3.270 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.765 4.460 2.150 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.500 -0.235 13.440 0.235 ;
        RECT  12.160 -0.235 12.500 0.465 ;
        RECT  11.235 -0.235 12.160 0.235 ;
        RECT  10.895 -0.235 11.235 0.760 ;
        RECT  8.275 -0.235 10.895 0.235 ;
        RECT  7.935 -0.235 8.275 0.730 ;
        RECT  4.675 -0.235 7.935 0.235 ;
        RECT  4.335 -0.235 4.675 0.465 ;
        RECT  3.660 -0.235 4.335 0.235 ;
        RECT  3.320 -0.235 3.660 0.465 ;
        RECT  1.240 -0.235 3.320 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.500 3.685 13.440 4.155 ;
        RECT  12.160 3.310 12.500 4.155 ;
        RECT  11.275 3.685 12.160 4.155 ;
        RECT  10.935 3.310 11.275 4.155 ;
        RECT  8.285 3.685 10.935 4.155 ;
        RECT  7.925 3.190 8.285 4.155 ;
        RECT  4.720 3.685 7.925 4.155 ;
        RECT  4.380 3.455 4.720 4.155 ;
        RECT  3.660 3.685 4.380 4.155 ;
        RECT  3.320 3.455 3.660 4.155 ;
        RECT  1.240 3.685 3.320 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.200 1.600 12.725 1.940 ;
        RECT  11.970 0.990 12.200 2.750 ;
        RECT  11.100 0.990 11.970 1.220 ;
        RECT  11.655 2.520 11.970 2.750 ;
        RECT  11.485 1.565 11.715 2.290 ;
        RECT  11.205 2.060 11.485 2.290 ;
        RECT  10.975 2.060 11.205 2.995 ;
        RECT  10.870 0.990 11.100 1.830 ;
        RECT  9.700 2.765 10.975 2.995 ;
        RECT  10.530 1.600 10.870 1.830 ;
        RECT  10.300 2.300 10.535 2.530 ;
        RECT  10.300 0.990 10.475 1.220 ;
        RECT  8.990 3.225 10.305 3.455 ;
        RECT  10.070 0.990 10.300 2.530 ;
        RECT  9.470 0.910 9.700 2.995 ;
        RECT  9.010 0.960 9.240 2.500 ;
        RECT  7.940 0.960 9.010 1.190 ;
        RECT  8.695 2.270 9.010 2.500 ;
        RECT  8.760 2.730 8.990 3.455 ;
        RECT  7.515 2.730 8.760 2.960 ;
        RECT  8.435 1.560 8.740 1.900 ;
        RECT  8.205 1.560 8.435 2.415 ;
        RECT  7.030 2.185 8.205 2.415 ;
        RECT  7.710 0.960 7.940 1.890 ;
        RECT  7.285 2.730 7.515 3.375 ;
        RECT  5.610 3.145 7.285 3.375 ;
        RECT  6.850 0.935 7.030 2.415 ;
        RECT  6.800 0.935 6.850 2.905 ;
        RECT  6.620 2.185 6.800 2.905 ;
        RECT  6.080 0.465 6.310 2.850 ;
        RECT  5.135 0.465 6.080 0.695 ;
        RECT  5.845 2.620 6.080 2.850 ;
        RECT  5.610 1.615 5.845 1.955 ;
        RECT  5.380 0.925 5.610 3.375 ;
        RECT  5.375 2.505 5.380 3.375 ;
        RECT  5.195 2.505 5.375 2.845 ;
        RECT  4.905 0.465 5.135 0.925 ;
        RECT  4.965 1.750 5.130 2.090 ;
        RECT  4.735 1.155 4.965 2.790 ;
        RECT  2.640 0.695 4.905 0.925 ;
        RECT  3.920 1.155 4.735 1.385 ;
        RECT  3.820 2.560 4.735 2.790 ;
        RECT  2.415 0.695 2.640 2.780 ;
        RECT  2.410 0.695 2.415 3.355 ;
        RECT  2.130 0.695 2.410 0.925 ;
        RECT  2.185 2.545 2.410 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFQD0BWP7T

MACRO SDFQD1BWP7T
    CLASS CORE ;
    FOREIGN SDFQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.1850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.530 0.470 13.860 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.470 1.760 4.620 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.005 -0.235 14.000 0.235 ;
        RECT  12.775 -0.235 13.005 1.255 ;
        RECT  11.625 -0.235 12.775 0.235 ;
        RECT  11.285 -0.235 11.625 0.670 ;
        RECT  8.510 -0.235 11.285 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.900 -0.235 4.575 0.235 ;
        RECT  3.560 -0.235 3.900 0.465 ;
        RECT  1.240 -0.235 3.560 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.005 3.685 14.000 4.155 ;
        RECT  12.775 2.255 13.005 4.155 ;
        RECT  11.635 3.685 12.775 4.155 ;
        RECT  11.295 3.250 11.635 4.155 ;
        RECT  8.520 3.685 11.295 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.960 3.685 8.160 4.155 ;
        RECT  4.620 3.455 4.960 4.155 ;
        RECT  3.780 3.685 4.620 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.240 3.685 3.440 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.545 1.600 13.265 1.940 ;
        RECT  12.315 1.020 12.545 2.795 ;
        RECT  12.300 1.020 12.315 1.250 ;
        RECT  12.300 2.565 12.315 2.795 ;
        RECT  12.070 0.495 12.300 1.250 ;
        RECT  12.070 2.565 12.300 3.380 ;
        RECT  11.845 1.565 12.075 2.310 ;
        RECT  11.465 1.020 12.070 1.250 ;
        RECT  11.565 2.080 11.845 2.310 ;
        RECT  11.335 2.080 11.565 2.995 ;
        RECT  11.235 1.020 11.465 1.830 ;
        RECT  9.975 2.765 11.335 2.995 ;
        RECT  10.850 1.600 11.235 1.830 ;
        RECT  10.535 2.300 10.830 2.530 ;
        RECT  10.535 0.990 10.790 1.220 ;
        RECT  9.225 3.225 10.540 3.455 ;
        RECT  10.305 0.990 10.535 2.530 ;
        RECT  9.745 0.910 9.975 2.995 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.375 ;
        RECT  5.845 3.145 7.520 3.375 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.615 6.080 1.955 ;
        RECT  5.615 0.925 5.845 3.375 ;
        RECT  5.375 2.560 5.615 2.790 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.090 ;
        RECT  2.600 0.695 5.145 0.925 ;
        RECT  4.240 1.155 5.140 1.385 ;
        RECT  4.240 2.505 4.345 2.845 ;
        RECT  4.010 1.155 4.240 2.845 ;
        RECT  2.445 0.695 2.600 2.780 ;
        RECT  2.370 0.695 2.445 3.355 ;
        RECT  2.195 0.695 2.370 0.925 ;
        RECT  2.215 2.545 2.370 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFQD1BWP7T

MACRO SDFQD2BWP7T
    CLASS CORE ;
    FOREIGN SDFQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.605 1.045 13.860 2.730 ;
        RECT  13.580 0.465 13.605 3.310 ;
        RECT  13.375 0.465 13.580 1.280 ;
        RECT  13.375 2.500 13.580 3.310 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.470 1.760 4.620 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 -0.235 14.560 0.235 ;
        RECT  14.095 -0.235 14.325 1.230 ;
        RECT  12.885 -0.235 14.095 0.235 ;
        RECT  12.655 -0.235 12.885 1.255 ;
        RECT  11.420 -0.235 12.655 0.235 ;
        RECT  11.080 -0.235 11.420 0.745 ;
        RECT  8.510 -0.235 11.080 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.900 -0.235 4.575 0.235 ;
        RECT  3.560 -0.235 3.900 0.465 ;
        RECT  1.240 -0.235 3.560 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 3.685 14.560 4.155 ;
        RECT  14.095 2.255 14.325 4.155 ;
        RECT  12.885 3.685 14.095 4.155 ;
        RECT  12.655 2.255 12.885 4.155 ;
        RECT  11.450 3.685 12.655 4.155 ;
        RECT  11.110 2.545 11.450 4.155 ;
        RECT  8.520 3.685 11.110 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.960 3.685 8.160 4.155 ;
        RECT  4.620 3.455 4.960 4.155 ;
        RECT  3.780 3.685 4.620 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.240 3.685 3.440 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.420 1.600 13.265 1.940 ;
        RECT  12.190 1.020 12.420 2.795 ;
        RECT  12.165 1.020 12.190 1.250 ;
        RECT  12.165 2.565 12.190 2.795 ;
        RECT  11.935 0.495 12.165 1.250 ;
        RECT  11.935 2.565 12.165 3.380 ;
        RECT  11.710 1.590 11.940 2.310 ;
        RECT  11.280 1.020 11.935 1.250 ;
        RECT  9.975 2.080 11.710 2.310 ;
        RECT  11.050 1.020 11.280 1.830 ;
        RECT  10.675 1.600 11.050 1.830 ;
        RECT  9.225 3.225 10.425 3.455 ;
        RECT  9.745 0.910 9.975 2.850 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.375 ;
        RECT  5.845 3.145 7.520 3.375 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.615 6.080 1.955 ;
        RECT  5.615 0.925 5.845 3.375 ;
        RECT  5.375 2.560 5.615 2.790 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.090 ;
        RECT  2.600 0.695 5.145 0.925 ;
        RECT  4.240 1.155 5.140 1.385 ;
        RECT  4.240 2.505 4.345 2.845 ;
        RECT  4.010 1.155 4.240 2.845 ;
        RECT  2.445 0.695 2.600 2.780 ;
        RECT  2.370 0.695 2.445 3.355 ;
        RECT  2.195 0.695 2.370 0.925 ;
        RECT  2.215 2.545 2.370 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFQD2BWP7T

MACRO SDFQND0BWP7T
    CLASS CORE ;
    FOREIGN SDFQND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5925 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.530 0.505 13.860 3.375 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.470 1.760 4.620 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.080 -0.235 14.000 0.235 ;
        RECT  12.740 -0.235 13.080 0.800 ;
        RECT  11.605 -0.235 12.740 0.235 ;
        RECT  11.375 -0.235 11.605 0.765 ;
        RECT  8.510 -0.235 11.375 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.900 -0.235 4.575 0.235 ;
        RECT  3.560 -0.235 3.900 0.465 ;
        RECT  1.240 -0.235 3.560 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.060 3.685 14.000 4.155 ;
        RECT  12.720 3.250 13.060 4.155 ;
        RECT  11.635 3.685 12.720 4.155 ;
        RECT  11.295 3.290 11.635 4.155 ;
        RECT  8.520 3.685 11.295 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.960 3.685 8.160 4.155 ;
        RECT  4.620 3.455 4.960 4.155 ;
        RECT  3.780 3.685 4.620 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.240 3.685 3.440 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.960 1.590 13.190 3.020 ;
        RECT  10.865 2.790 12.960 3.020 ;
        RECT  12.405 1.075 12.635 2.560 ;
        RECT  12.325 1.075 12.405 1.310 ;
        RECT  11.340 2.330 12.405 2.560 ;
        RECT  12.095 0.465 12.325 1.310 ;
        RECT  11.850 1.650 12.130 1.880 ;
        RECT  11.620 1.095 11.850 1.880 ;
        RECT  11.145 1.095 11.620 1.325 ;
        RECT  11.110 1.630 11.340 2.560 ;
        RECT  10.915 0.465 11.145 1.325 ;
        RECT  10.850 1.630 11.110 1.860 ;
        RECT  9.965 0.465 10.915 0.695 ;
        RECT  10.635 2.300 10.865 3.020 ;
        RECT  10.535 0.935 10.685 1.275 ;
        RECT  10.535 2.300 10.635 2.530 ;
        RECT  10.305 0.935 10.535 2.530 ;
        RECT  9.225 3.225 10.530 3.455 ;
        RECT  9.735 0.465 9.965 2.850 ;
        RECT  9.245 0.960 9.475 2.500 ;
        RECT  8.175 0.960 9.245 1.190 ;
        RECT  8.930 2.270 9.245 2.500 ;
        RECT  8.995 2.730 9.225 3.455 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.670 1.560 8.975 1.900 ;
        RECT  8.440 1.560 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.375 ;
        RECT  5.845 3.145 7.520 3.375 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.615 6.080 1.955 ;
        RECT  5.615 0.925 5.845 3.375 ;
        RECT  5.375 2.560 5.615 2.790 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.090 ;
        RECT  2.600 0.695 5.145 0.925 ;
        RECT  4.240 1.155 5.140 1.385 ;
        RECT  4.240 2.505 4.345 2.845 ;
        RECT  4.010 1.155 4.240 2.845 ;
        RECT  2.445 0.695 2.600 2.780 ;
        RECT  2.370 0.695 2.445 3.355 ;
        RECT  2.195 0.695 2.370 0.925 ;
        RECT  2.215 2.545 2.370 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFQND0BWP7T

MACRO SDFQND1BWP7T
    CLASS CORE ;
    FOREIGN SDFQND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.000 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5013 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.530 0.470 13.860 3.310 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.3924 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 1.725 3.780 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.760 4.900 2.710 ;
        RECT  4.470 1.760 4.620 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.025 -0.235 14.000 0.235 ;
        RECT  12.795 -0.235 13.025 1.255 ;
        RECT  11.605 -0.235 12.795 0.235 ;
        RECT  11.375 -0.235 11.605 0.725 ;
        RECT  8.510 -0.235 11.375 0.235 ;
        RECT  8.170 -0.235 8.510 0.730 ;
        RECT  4.915 -0.235 8.170 0.235 ;
        RECT  4.575 -0.235 4.915 0.465 ;
        RECT  3.900 -0.235 4.575 0.235 ;
        RECT  3.560 -0.235 3.900 0.465 ;
        RECT  1.240 -0.235 3.560 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.060 3.685 14.000 4.155 ;
        RECT  12.720 3.250 13.060 4.155 ;
        RECT  11.585 3.685 12.720 4.155 ;
        RECT  11.245 3.250 11.585 4.155 ;
        RECT  8.520 3.685 11.245 4.155 ;
        RECT  8.160 3.190 8.520 4.155 ;
        RECT  4.960 3.685 8.160 4.155 ;
        RECT  4.620 3.455 4.960 4.155 ;
        RECT  3.780 3.685 4.620 4.155 ;
        RECT  3.440 3.455 3.780 4.155 ;
        RECT  1.240 3.685 3.440 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.935 1.590 13.165 3.020 ;
        RECT  10.930 2.790 12.935 3.020 ;
        RECT  12.315 0.465 12.545 2.560 ;
        RECT  12.095 0.465 12.315 0.805 ;
        RECT  11.390 2.330 12.315 2.560 ;
        RECT  11.850 1.595 12.075 1.945 ;
        RECT  11.620 0.975 11.850 1.945 ;
        RECT  11.145 0.975 11.620 1.205 ;
        RECT  11.160 1.630 11.390 2.560 ;
        RECT  10.850 1.630 11.160 1.860 ;
        RECT  10.915 0.465 11.145 1.205 ;
        RECT  10.700 2.300 10.930 3.020 ;
        RECT  9.965 0.465 10.915 0.695 ;
        RECT  10.535 2.300 10.700 2.530 ;
        RECT  10.535 0.935 10.685 1.275 ;
        RECT  10.305 0.935 10.535 2.530 ;
        RECT  9.225 3.125 10.430 3.355 ;
        RECT  9.735 0.465 9.965 2.850 ;
        RECT  9.265 0.960 9.495 2.500 ;
        RECT  8.175 0.960 9.265 1.190 ;
        RECT  8.930 2.270 9.265 2.500 ;
        RECT  8.995 2.730 9.225 3.355 ;
        RECT  8.670 1.615 9.030 1.845 ;
        RECT  7.750 2.730 8.995 2.960 ;
        RECT  8.440 1.615 8.670 2.415 ;
        RECT  7.265 2.185 8.440 2.415 ;
        RECT  7.945 0.960 8.175 1.890 ;
        RECT  7.520 2.730 7.750 3.375 ;
        RECT  5.845 3.145 7.520 3.375 ;
        RECT  7.085 0.935 7.265 2.415 ;
        RECT  7.035 0.935 7.085 2.905 ;
        RECT  6.855 2.185 7.035 2.905 ;
        RECT  6.315 0.465 6.545 2.850 ;
        RECT  5.375 0.465 6.315 0.695 ;
        RECT  6.080 2.620 6.315 2.850 ;
        RECT  5.845 1.615 6.080 1.955 ;
        RECT  5.615 0.925 5.845 3.375 ;
        RECT  5.375 2.560 5.615 2.790 ;
        RECT  5.145 0.465 5.375 0.925 ;
        RECT  5.140 1.155 5.370 2.090 ;
        RECT  2.600 0.695 5.145 0.925 ;
        RECT  4.240 1.155 5.140 1.385 ;
        RECT  4.240 2.505 4.345 2.845 ;
        RECT  4.010 1.155 4.240 2.845 ;
        RECT  2.445 0.695 2.600 2.780 ;
        RECT  2.370 0.695 2.445 3.355 ;
        RECT  2.195 0.695 2.370 0.925 ;
        RECT  2.215 2.545 2.370 3.355 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFQND1BWP7T

MACRO SDFQND2BWP7T
    CLASS CORE ;
    FOREIGN SDFQND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.560 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.5094 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.605 1.065 13.860 2.730 ;
        RECT  13.580 0.470 13.605 3.310 ;
        RECT  13.375 0.470 13.580 1.295 ;
        RECT  13.375 2.500 13.580 3.310 ;
        END
    END QN
    PIN D
        ANTENNAGATEAREA 0.4005 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.725 3.310 2.160 ;
        RECT  2.940 1.725 3.220 2.710 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 1.760 4.520 2.150 ;
        RECT  3.575 1.210 3.805 2.150 ;
        RECT  3.500 1.210 3.575 1.590 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 -0.235 14.560 0.235 ;
        RECT  14.095 -0.235 14.325 1.230 ;
        RECT  12.885 -0.235 14.095 0.235 ;
        RECT  12.655 -0.235 12.885 1.255 ;
        RECT  11.465 -0.235 12.655 0.235 ;
        RECT  11.235 -0.235 11.465 0.725 ;
        RECT  8.370 -0.235 11.235 0.235 ;
        RECT  8.030 -0.235 8.370 0.730 ;
        RECT  4.775 -0.235 8.030 0.235 ;
        RECT  4.435 -0.235 4.775 0.465 ;
        RECT  3.805 -0.235 4.435 0.235 ;
        RECT  3.465 -0.235 3.805 0.465 ;
        RECT  1.240 -0.235 3.465 0.235 ;
        RECT  0.900 -0.235 1.240 0.870 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.325 3.685 14.560 4.155 ;
        RECT  14.095 2.250 14.325 4.155 ;
        RECT  12.940 3.685 14.095 4.155 ;
        RECT  12.600 3.250 12.940 4.155 ;
        RECT  11.445 3.685 12.600 4.155 ;
        RECT  11.105 3.250 11.445 4.155 ;
        RECT  8.380 3.685 11.105 4.155 ;
        RECT  8.020 3.190 8.380 4.155 ;
        RECT  4.820 3.685 8.020 4.155 ;
        RECT  4.480 3.455 4.820 4.155 ;
        RECT  3.645 3.685 4.480 4.155 ;
        RECT  3.305 3.455 3.645 4.155 ;
        RECT  1.240 3.685 3.305 4.155 ;
        RECT  0.900 2.940 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.795 1.590 13.025 3.020 ;
        RECT  10.790 2.790 12.795 3.020 ;
        RECT  12.185 1.075 12.405 2.560 ;
        RECT  12.175 0.495 12.185 2.560 ;
        RECT  11.955 0.495 12.175 1.310 ;
        RECT  11.250 2.330 12.175 2.560 ;
        RECT  11.710 1.595 11.935 1.945 ;
        RECT  11.480 0.975 11.710 1.945 ;
        RECT  11.005 0.975 11.480 1.205 ;
        RECT  11.020 1.630 11.250 2.560 ;
        RECT  10.710 1.630 11.020 1.860 ;
        RECT  10.775 0.465 11.005 1.205 ;
        RECT  10.560 2.300 10.790 3.020 ;
        RECT  9.825 0.465 10.775 0.695 ;
        RECT  10.395 2.300 10.560 2.530 ;
        RECT  10.395 0.935 10.545 1.275 ;
        RECT  10.165 0.935 10.395 2.530 ;
        RECT  9.085 3.125 10.290 3.355 ;
        RECT  9.595 0.465 9.825 2.850 ;
        RECT  9.125 0.960 9.355 2.500 ;
        RECT  8.035 0.960 9.125 1.190 ;
        RECT  8.790 2.270 9.125 2.500 ;
        RECT  8.855 2.730 9.085 3.355 ;
        RECT  8.530 1.615 8.890 1.845 ;
        RECT  7.610 2.730 8.855 2.960 ;
        RECT  8.300 1.615 8.530 2.415 ;
        RECT  7.125 2.185 8.300 2.415 ;
        RECT  7.805 0.960 8.035 1.890 ;
        RECT  7.380 2.730 7.610 3.375 ;
        RECT  5.705 3.145 7.380 3.375 ;
        RECT  6.945 0.935 7.125 2.415 ;
        RECT  6.895 0.935 6.945 2.905 ;
        RECT  6.715 2.185 6.895 2.905 ;
        RECT  6.175 0.465 6.405 2.850 ;
        RECT  5.235 0.465 6.175 0.695 ;
        RECT  5.940 2.620 6.175 2.850 ;
        RECT  5.705 1.615 5.940 1.955 ;
        RECT  5.475 0.925 5.705 3.375 ;
        RECT  5.295 2.505 5.475 2.850 ;
        RECT  5.025 1.750 5.245 2.090 ;
        RECT  5.005 0.465 5.235 0.925 ;
        RECT  4.795 1.155 5.025 2.790 ;
        RECT  2.640 0.695 5.005 0.925 ;
        RECT  4.050 1.155 4.795 1.385 ;
        RECT  3.920 2.560 4.795 2.790 ;
        RECT  2.410 0.695 2.640 3.055 ;
        RECT  2.130 0.695 2.410 0.925 ;
        RECT  2.090 2.815 2.410 3.055 ;
        RECT  2.000 1.725 2.135 2.065 ;
        RECT  1.770 1.130 2.000 2.065 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFQND2BWP7T

MACRO SDFSND0BWP7T
    CLASS CORE ;
    FOREIGN SDFSND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.715 2.940 12.055 3.370 ;
        RECT  10.485 2.940 11.715 3.220 ;
        RECT  10.255 2.730 10.485 3.220 ;
        RECT  8.730 2.730 10.255 2.960 ;
        RECT  8.500 2.730 8.730 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.565 16.660 2.720 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.120 15.540 2.660 ;
        RECT  15.125 1.120 15.260 1.350 ;
        RECT  14.840 2.430 15.260 2.660 ;
        RECT  14.895 0.560 15.125 1.350 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.380 1.605 3.500 1.945 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.630 4.900 2.710 ;
        RECT  4.485 1.630 4.620 1.970 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.860 ;
        RECT  13.565 -0.235 15.560 0.235 ;
        RECT  13.225 -0.235 13.565 0.860 ;
        RECT  8.530 -0.235 13.225 0.235 ;
        RECT  8.190 -0.235 8.530 0.960 ;
        RECT  4.135 -0.235 8.190 0.235 ;
        RECT  3.795 -0.235 4.135 0.465 ;
        RECT  1.240 -0.235 3.795 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.830 3.685 16.800 4.155 ;
        RECT  15.490 3.455 15.830 4.155 ;
        RECT  13.715 3.685 15.490 4.155 ;
        RECT  13.375 3.455 13.715 4.155 ;
        RECT  12.690 3.685 13.375 4.155 ;
        RECT  12.350 3.450 12.690 4.155 ;
        RECT  9.920 3.685 12.350 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.975 3.685 7.980 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.410 16.085 3.225 ;
        RECT  13.325 2.995 15.855 3.225 ;
        RECT  14.610 1.635 15.030 1.865 ;
        RECT  14.425 0.630 14.610 2.230 ;
        RECT  14.380 0.630 14.425 2.725 ;
        RECT  13.990 0.630 14.380 0.860 ;
        RECT  14.195 2.000 14.380 2.725 ;
        RECT  13.080 2.000 14.195 2.230 ;
        RECT  13.805 1.205 14.035 1.750 ;
        RECT  12.800 1.205 13.805 1.435 ;
        RECT  13.090 2.465 13.325 3.225 ;
        RECT  11.845 2.465 13.090 2.695 ;
        RECT  12.740 1.780 13.080 2.230 ;
        RECT  12.570 0.465 12.800 1.435 ;
        RECT  10.580 0.465 12.570 0.695 ;
        RECT  11.845 0.990 12.170 1.220 ;
        RECT  11.615 0.990 11.845 2.695 ;
        RECT  11.015 0.990 11.615 1.220 ;
        RECT  10.895 1.615 11.125 2.585 ;
        RECT  10.580 1.615 10.895 1.845 ;
        RECT  10.350 0.465 10.580 1.845 ;
        RECT  10.030 2.270 10.460 2.500 ;
        RECT  9.800 0.935 10.030 2.500 ;
        RECT  9.510 0.935 9.800 1.165 ;
        RECT  8.195 2.270 9.800 2.500 ;
        RECT  8.965 1.640 9.490 1.870 ;
        RECT  8.735 1.190 8.965 1.870 ;
        RECT  7.240 1.190 8.735 1.420 ;
        RECT  7.965 1.655 8.195 2.500 ;
        RECT  7.100 0.660 7.240 1.420 ;
        RECT  7.010 0.660 7.100 3.085 ;
        RECT  6.870 1.190 7.010 3.085 ;
        RECT  6.380 0.705 6.600 2.505 ;
        RECT  6.370 0.705 6.380 3.225 ;
        RECT  6.235 0.705 6.370 0.935 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.880 1.505 6.095 1.845 ;
        RECT  5.650 0.910 5.880 2.765 ;
        RECT  5.590 0.910 5.650 1.270 ;
        RECT  5.390 2.535 5.650 2.765 ;
        RECT  5.360 1.620 5.385 1.960 ;
        RECT  5.130 0.980 5.360 1.960 ;
        RECT  4.255 0.980 5.130 1.210 ;
        RECT  4.255 2.420 4.360 2.760 ;
        RECT  4.025 0.980 4.255 2.760 ;
        RECT  3.315 2.995 3.545 3.450 ;
        RECT  2.600 3.220 3.315 3.450 ;
        RECT  3.095 0.465 3.200 1.275 ;
        RECT  2.970 0.465 3.095 2.925 ;
        RECT  2.865 1.080 2.970 2.925 ;
        RECT  2.480 1.085 2.600 3.450 ;
        RECT  2.370 0.465 2.480 3.450 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFSND0BWP7T

MACRO SDFSND1BWP7T
    CLASS CORE ;
    FOREIGN SDFSND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.800 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.715 2.940 12.055 3.340 ;
        RECT  10.485 2.940 11.715 3.220 ;
        RECT  10.255 2.730 10.485 3.220 ;
        RECT  8.730 2.730 10.255 2.960 ;
        RECT  8.500 2.730 8.730 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.330 0.470 16.660 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.260 1.075 15.540 2.560 ;
        RECT  15.125 1.075 15.260 1.305 ;
        RECT  14.840 2.330 15.260 2.560 ;
        RECT  14.895 0.465 15.125 1.305 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.380 1.605 3.500 1.945 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.630 4.900 2.710 ;
        RECT  4.485 1.630 4.620 1.970 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 -0.235 16.800 0.235 ;
        RECT  15.560 -0.235 15.900 0.810 ;
        RECT  13.570 -0.235 15.560 0.235 ;
        RECT  13.230 -0.235 13.570 0.930 ;
        RECT  8.530 -0.235 13.230 0.235 ;
        RECT  8.190 -0.235 8.530 0.960 ;
        RECT  4.135 -0.235 8.190 0.235 ;
        RECT  3.795 -0.235 4.135 0.465 ;
        RECT  1.240 -0.235 3.795 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.900 3.685 16.800 4.155 ;
        RECT  15.560 3.250 15.900 4.155 ;
        RECT  13.715 3.685 15.560 4.155 ;
        RECT  13.375 3.455 13.715 4.155 ;
        RECT  12.690 3.685 13.375 4.155 ;
        RECT  12.350 3.450 12.690 4.155 ;
        RECT  9.920 3.685 12.350 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.975 3.685 7.980 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.855 1.600 16.085 3.020 ;
        RECT  15.085 2.790 15.855 3.020 ;
        RECT  14.855 2.790 15.085 3.225 ;
        RECT  14.610 1.635 15.030 1.865 ;
        RECT  13.325 2.995 14.855 3.225 ;
        RECT  14.425 0.680 14.610 2.230 ;
        RECT  14.380 0.680 14.425 2.765 ;
        RECT  13.990 0.680 14.380 0.910 ;
        RECT  14.195 2.000 14.380 2.765 ;
        RECT  13.080 2.000 14.195 2.230 ;
        RECT  13.745 1.205 14.090 1.770 ;
        RECT  12.800 1.205 13.745 1.435 ;
        RECT  13.090 2.465 13.325 3.225 ;
        RECT  11.845 2.465 13.090 2.695 ;
        RECT  12.740 1.780 13.080 2.230 ;
        RECT  12.570 0.465 12.800 1.435 ;
        RECT  10.580 0.465 12.570 0.695 ;
        RECT  11.845 0.990 12.170 1.220 ;
        RECT  11.615 0.990 11.845 2.695 ;
        RECT  11.015 0.990 11.615 1.220 ;
        RECT  10.895 1.615 11.125 2.585 ;
        RECT  10.580 1.615 10.895 1.845 ;
        RECT  10.350 0.465 10.580 1.845 ;
        RECT  10.030 2.270 10.460 2.500 ;
        RECT  9.800 0.935 10.030 2.500 ;
        RECT  9.510 0.935 9.800 1.165 ;
        RECT  8.195 2.270 9.800 2.500 ;
        RECT  8.965 1.640 9.490 1.870 ;
        RECT  8.735 1.190 8.965 1.870 ;
        RECT  7.240 1.190 8.735 1.420 ;
        RECT  7.965 1.655 8.195 2.500 ;
        RECT  7.100 0.660 7.240 1.420 ;
        RECT  7.010 0.660 7.100 3.085 ;
        RECT  6.870 1.190 7.010 3.085 ;
        RECT  6.380 0.705 6.600 2.505 ;
        RECT  6.370 0.705 6.380 3.225 ;
        RECT  6.235 0.705 6.370 0.935 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.880 1.505 6.095 1.845 ;
        RECT  5.650 0.910 5.880 2.765 ;
        RECT  5.590 0.910 5.650 1.270 ;
        RECT  5.390 2.535 5.650 2.765 ;
        RECT  5.360 1.620 5.385 1.960 ;
        RECT  5.130 0.980 5.360 1.960 ;
        RECT  4.255 0.980 5.130 1.210 ;
        RECT  4.255 2.420 4.360 2.760 ;
        RECT  4.025 0.980 4.255 2.760 ;
        RECT  3.315 2.995 3.545 3.450 ;
        RECT  2.600 3.220 3.315 3.450 ;
        RECT  3.095 0.465 3.200 1.275 ;
        RECT  2.970 0.465 3.095 2.925 ;
        RECT  2.865 1.080 2.970 2.925 ;
        RECT  2.480 1.085 2.600 3.450 ;
        RECT  2.370 0.465 2.480 3.450 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFSND1BWP7T

MACRO SDFSND2BWP7T
    CLASS CORE ;
    FOREIGN SDFSND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.4761 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.715 2.940 12.055 3.370 ;
        RECT  10.485 2.940 11.715 3.220 ;
        RECT  10.255 2.730 10.485 3.220 ;
        RECT  8.730 2.730 10.255 2.960 ;
        RECT  8.500 2.730 8.730 3.155 ;
        END
    END SDN
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 1.055 17.220 2.690 ;
        RECT  16.940 0.465 16.965 3.310 ;
        RECT  16.730 0.465 16.940 1.285 ;
        RECT  16.735 2.460 16.940 3.310 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.240 0.465 15.585 2.560 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.380 1.605 3.500 1.945 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.630 4.900 2.710 ;
        RECT  4.485 1.630 4.620 1.970 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 -0.235 17.920 0.235 ;
        RECT  17.455 -0.235 17.685 1.245 ;
        RECT  16.300 -0.235 17.455 0.235 ;
        RECT  15.960 -0.235 16.300 1.180 ;
        RECT  14.820 -0.235 15.960 0.235 ;
        RECT  14.480 -0.235 14.820 0.480 ;
        RECT  13.360 -0.235 14.480 0.235 ;
        RECT  13.020 -0.235 13.360 0.910 ;
        RECT  8.530 -0.235 13.020 0.235 ;
        RECT  8.190 -0.235 8.530 0.960 ;
        RECT  4.135 -0.235 8.190 0.235 ;
        RECT  3.795 -0.235 4.135 0.465 ;
        RECT  1.240 -0.235 3.795 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.685 3.685 17.920 4.155 ;
        RECT  17.455 2.255 17.685 4.155 ;
        RECT  16.300 3.685 17.455 4.155 ;
        RECT  15.960 3.250 16.300 4.155 ;
        RECT  14.860 3.685 15.960 4.155 ;
        RECT  14.520 3.250 14.860 4.155 ;
        RECT  12.705 3.685 14.520 4.155 ;
        RECT  12.365 3.025 12.705 4.155 ;
        RECT  9.920 3.685 12.365 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.975 3.685 7.980 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.255 1.600 16.485 3.020 ;
        RECT  13.380 2.790 16.255 3.020 ;
        RECT  14.770 0.730 15.000 2.245 ;
        RECT  13.720 0.730 14.770 0.960 ;
        RECT  14.140 2.015 14.770 2.245 ;
        RECT  14.030 1.215 14.375 1.785 ;
        RECT  13.800 2.015 14.140 2.560 ;
        RECT  12.745 1.215 14.030 1.445 ;
        RECT  13.130 2.015 13.800 2.245 ;
        RECT  13.150 2.475 13.380 3.315 ;
        RECT  11.845 2.475 13.150 2.705 ;
        RECT  12.785 1.675 13.130 2.245 ;
        RECT  12.515 0.465 12.745 1.445 ;
        RECT  10.580 0.465 12.515 0.695 ;
        RECT  11.845 0.990 12.155 1.220 ;
        RECT  11.615 0.990 11.845 2.705 ;
        RECT  11.015 0.990 11.615 1.220 ;
        RECT  10.895 1.615 11.125 2.585 ;
        RECT  10.580 1.615 10.895 1.845 ;
        RECT  10.350 0.465 10.580 1.845 ;
        RECT  10.030 2.270 10.460 2.500 ;
        RECT  9.800 0.935 10.030 2.500 ;
        RECT  9.510 0.935 9.800 1.165 ;
        RECT  8.195 2.270 9.800 2.500 ;
        RECT  8.965 1.640 9.490 1.870 ;
        RECT  8.735 1.190 8.965 1.870 ;
        RECT  7.240 1.190 8.735 1.420 ;
        RECT  7.965 1.655 8.195 2.500 ;
        RECT  7.100 0.660 7.240 1.420 ;
        RECT  7.010 0.660 7.100 3.085 ;
        RECT  6.870 1.190 7.010 3.085 ;
        RECT  6.380 0.705 6.600 2.505 ;
        RECT  6.370 0.705 6.380 3.225 ;
        RECT  6.235 0.705 6.370 0.935 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.880 1.505 6.095 1.845 ;
        RECT  5.650 0.910 5.880 2.765 ;
        RECT  5.590 0.910 5.650 1.270 ;
        RECT  5.390 2.535 5.650 2.765 ;
        RECT  5.360 1.620 5.385 1.960 ;
        RECT  5.130 0.980 5.360 1.960 ;
        RECT  4.255 0.980 5.130 1.210 ;
        RECT  4.255 2.420 4.360 2.760 ;
        RECT  4.025 0.980 4.255 2.760 ;
        RECT  3.315 2.995 3.545 3.450 ;
        RECT  2.600 3.220 3.315 3.450 ;
        RECT  3.095 0.465 3.200 1.275 ;
        RECT  2.970 0.465 3.095 2.925 ;
        RECT  2.865 1.080 2.970 2.925 ;
        RECT  2.480 1.085 2.600 3.450 ;
        RECT  2.370 0.465 2.480 3.450 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFSND2BWP7T

MACRO SDFSNQD0BWP7T
    CLASS CORE ;
    FOREIGN SDFSNQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.715 2.940 12.055 3.315 ;
        RECT  10.485 2.940 11.715 3.220 ;
        RECT  10.255 2.730 10.485 3.220 ;
        RECT  8.785 2.730 10.255 2.960 ;
        RECT  8.440 2.730 8.785 3.025 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.775 0.600 16.100 3.200 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.595 3.780 2.710 ;
        RECT  3.380 1.595 3.500 1.935 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.675 4.900 2.710 ;
        RECT  4.485 1.675 4.620 2.025 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.340 -0.235 16.240 0.235 ;
        RECT  15.000 -0.235 15.340 0.900 ;
        RECT  13.760 -0.235 15.000 0.235 ;
        RECT  13.420 -0.235 13.760 0.830 ;
        RECT  8.525 -0.235 13.420 0.235 ;
        RECT  8.185 -0.235 8.525 0.960 ;
        RECT  4.185 -0.235 8.185 0.235 ;
        RECT  3.845 -0.235 4.185 0.465 ;
        RECT  1.240 -0.235 3.845 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.340 3.685 16.240 4.155 ;
        RECT  15.000 2.915 15.340 4.155 ;
        RECT  13.900 3.685 15.000 4.155 ;
        RECT  13.560 2.650 13.900 4.155 ;
        RECT  12.690 3.685 13.560 4.155 ;
        RECT  12.350 3.450 12.690 4.155 ;
        RECT  9.920 3.685 12.350 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.975 3.685 7.980 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.980 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.585 1.655 15.545 1.885 ;
        RECT  14.355 0.550 14.585 2.905 ;
        RECT  13.275 2.000 14.355 2.230 ;
        RECT  13.745 1.190 14.090 1.770 ;
        RECT  12.955 1.190 13.745 1.420 ;
        RECT  12.935 1.780 13.275 2.230 ;
        RECT  12.875 2.465 13.105 2.940 ;
        RECT  12.725 0.465 12.955 1.420 ;
        RECT  11.845 2.465 12.875 2.695 ;
        RECT  10.580 0.465 12.725 0.695 ;
        RECT  11.845 0.990 12.305 1.220 ;
        RECT  11.615 0.990 11.845 2.695 ;
        RECT  11.015 0.990 11.615 1.220 ;
        RECT  10.895 1.615 11.125 2.585 ;
        RECT  10.580 1.615 10.895 1.845 ;
        RECT  10.350 0.465 10.580 1.845 ;
        RECT  10.070 2.270 10.460 2.500 ;
        RECT  9.840 0.930 10.070 2.500 ;
        RECT  9.490 0.930 9.840 1.160 ;
        RECT  8.190 2.270 9.840 2.500 ;
        RECT  8.965 1.645 9.555 1.875 ;
        RECT  8.735 1.190 8.965 1.875 ;
        RECT  7.240 1.190 8.735 1.420 ;
        RECT  7.960 1.650 8.190 2.500 ;
        RECT  7.100 0.660 7.240 1.420 ;
        RECT  7.010 0.660 7.100 3.085 ;
        RECT  6.870 1.190 7.010 3.085 ;
        RECT  6.380 0.705 6.600 2.505 ;
        RECT  6.370 0.705 6.380 3.225 ;
        RECT  6.235 0.705 6.370 0.935 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.880 1.505 6.095 1.845 ;
        RECT  5.650 0.920 5.880 2.765 ;
        RECT  5.590 0.920 5.650 1.260 ;
        RECT  5.390 2.535 5.650 2.765 ;
        RECT  5.360 1.660 5.390 2.000 ;
        RECT  5.130 0.975 5.360 2.000 ;
        RECT  4.240 0.975 5.130 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.450 ;
        RECT  2.600 3.220 3.315 3.450 ;
        RECT  3.095 0.465 3.200 1.275 ;
        RECT  2.970 0.465 3.095 2.855 ;
        RECT  2.865 1.080 2.970 2.855 ;
        RECT  2.480 1.085 2.600 3.450 ;
        RECT  2.370 0.465 2.480 3.450 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFSNQD0BWP7T

MACRO SDFSNQD1BWP7T
    CLASS CORE ;
    FOREIGN SDFSNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.3861 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.715 2.940 12.055 3.315 ;
        RECT  10.485 2.940 11.715 3.220 ;
        RECT  10.255 2.730 10.485 3.220 ;
        RECT  8.785 2.730 10.255 2.960 ;
        RECT  8.440 2.730 8.785 3.025 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.775 0.465 16.100 3.300 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.595 3.780 2.710 ;
        RECT  3.380 1.595 3.500 1.935 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.675 4.900 2.710 ;
        RECT  4.485 1.675 4.620 2.025 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.340 -0.235 16.240 0.235 ;
        RECT  15.000 -0.235 15.340 1.205 ;
        RECT  13.760 -0.235 15.000 0.235 ;
        RECT  13.420 -0.235 13.760 0.890 ;
        RECT  8.525 -0.235 13.420 0.235 ;
        RECT  8.185 -0.235 8.525 0.960 ;
        RECT  4.190 -0.235 8.185 0.235 ;
        RECT  3.850 -0.235 4.190 0.465 ;
        RECT  1.240 -0.235 3.850 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.340 3.685 16.240 4.155 ;
        RECT  15.000 2.555 15.340 4.155 ;
        RECT  13.920 3.685 15.000 4.155 ;
        RECT  13.580 2.540 13.920 4.155 ;
        RECT  12.690 3.685 13.580 4.155 ;
        RECT  12.350 3.450 12.690 4.155 ;
        RECT  9.920 3.685 12.350 4.155 ;
        RECT  9.580 3.190 9.920 4.155 ;
        RECT  8.210 3.685 9.580 4.155 ;
        RECT  7.980 3.130 8.210 4.155 ;
        RECT  4.975 3.685 7.980 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.980 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.585 1.655 15.545 1.885 ;
        RECT  14.355 0.465 14.585 3.315 ;
        RECT  13.275 2.000 14.355 2.230 ;
        RECT  13.745 1.190 14.090 1.770 ;
        RECT  12.955 1.190 13.745 1.420 ;
        RECT  12.935 1.780 13.275 2.230 ;
        RECT  11.845 2.465 13.170 2.695 ;
        RECT  12.725 0.465 12.955 1.420 ;
        RECT  10.580 0.465 12.725 0.695 ;
        RECT  11.845 0.990 12.305 1.220 ;
        RECT  11.615 0.990 11.845 2.695 ;
        RECT  11.015 0.990 11.615 1.220 ;
        RECT  10.895 1.615 11.125 2.585 ;
        RECT  10.580 1.615 10.895 1.845 ;
        RECT  10.350 0.465 10.580 1.845 ;
        RECT  10.070 2.270 10.460 2.500 ;
        RECT  9.840 0.930 10.070 2.500 ;
        RECT  9.485 0.930 9.840 1.160 ;
        RECT  8.190 2.270 9.840 2.500 ;
        RECT  8.965 1.635 9.555 1.865 ;
        RECT  8.735 1.190 8.965 1.865 ;
        RECT  7.240 1.190 8.735 1.420 ;
        RECT  7.960 1.650 8.190 2.500 ;
        RECT  7.100 0.660 7.240 1.420 ;
        RECT  7.010 0.660 7.100 3.085 ;
        RECT  6.870 1.190 7.010 3.085 ;
        RECT  6.380 0.705 6.600 2.505 ;
        RECT  6.370 0.705 6.380 3.225 ;
        RECT  6.235 0.705 6.370 0.935 ;
        RECT  6.150 2.275 6.370 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.880 1.505 6.095 1.845 ;
        RECT  5.650 0.920 5.880 2.765 ;
        RECT  5.590 0.920 5.650 1.260 ;
        RECT  5.390 2.535 5.650 2.765 ;
        RECT  5.360 1.660 5.390 2.000 ;
        RECT  5.130 0.975 5.360 2.000 ;
        RECT  4.240 0.975 5.130 1.205 ;
        RECT  4.240 2.425 4.360 2.765 ;
        RECT  4.010 0.975 4.240 2.765 ;
        RECT  3.315 2.995 3.545 3.450 ;
        RECT  2.600 3.220 3.315 3.450 ;
        RECT  3.095 0.465 3.200 1.275 ;
        RECT  2.970 0.465 3.095 2.855 ;
        RECT  2.865 1.080 2.970 2.855 ;
        RECT  2.480 1.085 2.600 3.450 ;
        RECT  2.370 0.465 2.480 3.450 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.935 0.520 3.165 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.165 ;
        RECT  0.115 1.130 0.235 3.165 ;
    END
END SDFSNQD1BWP7T

MACRO SDFSNQD2BWP7T
    CLASS CORE ;
    FOREIGN SDFSNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.240 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SE
    PIN SDN
        ANTENNAGATEAREA 0.3717 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.605 2.940 11.945 3.370 ;
        RECT  10.310 2.940 11.605 3.220 ;
        RECT  10.080 2.730 10.310 3.220 ;
        RECT  8.610 2.730 10.080 2.960 ;
        RECT  8.380 2.730 8.610 3.330 ;
        END
    END SDN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 1.100 15.540 2.675 ;
        RECT  15.260 0.465 15.285 3.335 ;
        RECT  15.055 0.465 15.260 1.355 ;
        RECT  15.055 2.360 15.260 3.335 ;
        END
    END Q
    PIN D
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.605 3.780 2.710 ;
        RECT  3.380 1.605 3.500 1.945 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.630 4.900 2.710 ;
        RECT  4.485 1.630 4.620 1.970 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 -0.235 16.240 0.235 ;
        RECT  15.775 -0.235 16.005 1.250 ;
        RECT  14.620 -0.235 15.775 0.235 ;
        RECT  14.280 -0.235 14.620 0.670 ;
        RECT  13.145 -0.235 14.280 0.235 ;
        RECT  12.915 -0.235 13.145 0.865 ;
        RECT  8.530 -0.235 12.915 0.235 ;
        RECT  8.190 -0.235 8.530 0.960 ;
        RECT  4.135 -0.235 8.190 0.235 ;
        RECT  3.795 -0.235 4.135 0.465 ;
        RECT  1.240 -0.235 3.795 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.005 3.685 16.240 4.155 ;
        RECT  15.775 2.245 16.005 4.155 ;
        RECT  14.620 3.685 15.775 4.155 ;
        RECT  14.280 3.250 14.620 4.155 ;
        RECT  12.525 3.685 14.280 4.155 ;
        RECT  12.185 2.995 12.525 4.155 ;
        RECT  9.785 3.685 12.185 4.155 ;
        RECT  9.445 3.190 9.785 4.155 ;
        RECT  8.050 3.685 9.445 4.155 ;
        RECT  7.820 3.130 8.050 4.155 ;
        RECT  4.975 3.685 7.820 4.155 ;
        RECT  4.635 3.455 4.975 4.155 ;
        RECT  4.115 3.685 4.635 4.155 ;
        RECT  3.775 3.455 4.115 4.155 ;
        RECT  1.240 3.685 3.775 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.530 1.075 14.760 2.245 ;
        RECT  13.845 1.075 14.530 1.305 ;
        RECT  13.900 2.015 14.530 2.245 ;
        RECT  13.385 1.555 14.135 1.785 ;
        RECT  13.560 2.015 13.900 2.610 ;
        RECT  13.615 0.885 13.845 1.305 ;
        RECT  12.815 2.015 13.560 2.245 ;
        RECT  13.155 1.215 13.385 1.785 ;
        RECT  13.060 3.060 13.245 3.290 ;
        RECT  12.555 1.215 13.155 1.445 ;
        RECT  12.830 2.475 13.060 3.290 ;
        RECT  11.710 2.475 12.830 2.705 ;
        RECT  12.575 1.705 12.815 2.245 ;
        RECT  12.325 0.465 12.555 1.445 ;
        RECT  10.385 0.465 12.325 0.695 ;
        RECT  11.710 0.990 11.960 1.250 ;
        RECT  11.480 0.990 11.710 2.705 ;
        RECT  10.820 0.990 11.480 1.220 ;
        RECT  10.760 1.615 10.990 2.585 ;
        RECT  10.385 1.615 10.760 1.845 ;
        RECT  10.155 0.465 10.385 1.845 ;
        RECT  9.885 2.270 10.285 2.500 ;
        RECT  9.655 0.935 9.885 2.500 ;
        RECT  9.375 0.935 9.655 1.165 ;
        RECT  8.010 2.270 9.655 2.500 ;
        RECT  9.195 1.585 9.425 1.935 ;
        RECT  8.965 1.585 9.195 1.815 ;
        RECT  8.735 1.190 8.965 1.815 ;
        RECT  7.240 1.190 8.735 1.420 ;
        RECT  7.780 1.875 8.010 2.500 ;
        RECT  7.100 0.855 7.240 1.420 ;
        RECT  7.010 0.855 7.100 2.735 ;
        RECT  6.870 1.190 7.010 2.735 ;
        RECT  6.380 0.705 6.600 2.310 ;
        RECT  6.370 0.705 6.380 3.225 ;
        RECT  6.235 0.705 6.370 0.935 ;
        RECT  6.150 2.080 6.370 3.225 ;
        RECT  3.545 2.995 6.150 3.225 ;
        RECT  5.880 1.505 6.095 1.845 ;
        RECT  5.650 0.910 5.880 2.765 ;
        RECT  5.590 0.910 5.650 1.270 ;
        RECT  5.390 2.535 5.650 2.765 ;
        RECT  5.360 1.620 5.385 1.960 ;
        RECT  5.130 0.980 5.360 1.960 ;
        RECT  4.255 0.980 5.130 1.210 ;
        RECT  4.255 2.420 4.360 2.760 ;
        RECT  4.025 0.980 4.255 2.760 ;
        RECT  3.315 2.995 3.545 3.450 ;
        RECT  2.600 3.220 3.315 3.450 ;
        RECT  3.095 0.465 3.200 1.275 ;
        RECT  2.970 0.465 3.095 2.925 ;
        RECT  2.865 1.080 2.970 2.925 ;
        RECT  2.480 1.085 2.600 3.450 ;
        RECT  2.370 0.465 2.480 3.450 ;
        RECT  2.250 0.465 2.370 1.290 ;
        RECT  2.090 2.820 2.370 3.050 ;
        RECT  2.000 1.810 2.135 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFSNQD2BWP7T

MACRO SDFXD0BWP7T
    CLASS CORE ;
    FOREIGN SDFXD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 1.750 7.160 2.150 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.750 6.020 2.150 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.5040 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.060 1.075 18.340 2.560 ;
        RECT  17.925 1.075 18.060 1.305 ;
        RECT  17.640 2.330 18.060 2.560 ;
        RECT  17.695 0.520 17.925 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.130 0.510 19.460 2.715 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4248 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.735 3.360 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2241 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.760 9.940 2.710 ;
        RECT  9.510 1.760 9.660 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.700 -0.235 19.600 0.235 ;
        RECT  18.360 -0.235 18.700 0.810 ;
        RECT  15.570 -0.235 18.360 0.235 ;
        RECT  15.230 -0.235 15.570 0.465 ;
        RECT  13.550 -0.235 15.230 0.235 ;
        RECT  13.210 -0.235 13.550 0.730 ;
        RECT  9.955 -0.235 13.210 0.235 ;
        RECT  9.615 -0.235 9.955 0.465 ;
        RECT  8.835 -0.235 9.615 0.235 ;
        RECT  8.495 -0.235 8.835 0.465 ;
        RECT  6.115 -0.235 8.495 0.235 ;
        RECT  5.775 -0.235 6.115 0.840 ;
        RECT  3.795 -0.235 5.775 0.235 ;
        RECT  3.455 -0.235 3.795 1.145 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.770 3.685 19.600 4.155 ;
        RECT  18.430 3.365 18.770 4.155 ;
        RECT  16.470 3.685 18.430 4.155 ;
        RECT  16.130 3.385 16.470 4.155 ;
        RECT  13.560 3.685 16.130 4.155 ;
        RECT  13.200 3.190 13.560 4.155 ;
        RECT  10.000 3.685 13.200 4.155 ;
        RECT  9.660 3.455 10.000 4.155 ;
        RECT  8.865 3.685 9.660 4.155 ;
        RECT  8.525 3.455 8.865 4.155 ;
        RECT  6.140 3.685 8.525 4.155 ;
        RECT  5.910 3.025 6.140 4.155 ;
        RECT  3.825 3.685 5.910 4.155 ;
        RECT  3.485 3.020 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.655 1.600 18.885 3.020 ;
        RECT  17.410 2.790 18.655 3.020 ;
        RECT  16.030 0.465 17.460 0.695 ;
        RECT  17.180 1.020 17.410 3.020 ;
        RECT  16.490 1.020 17.180 1.250 ;
        RECT  16.940 2.540 17.180 2.775 ;
        RECT  16.720 1.565 16.950 2.310 ;
        RECT  16.490 2.080 16.720 2.310 ;
        RECT  16.260 1.020 16.490 1.830 ;
        RECT  16.260 2.080 16.490 2.995 ;
        RECT  15.775 1.600 16.260 1.830 ;
        RECT  14.975 2.765 16.260 2.995 ;
        RECT  15.800 0.465 16.030 1.220 ;
        RECT  15.540 2.300 15.810 2.530 ;
        RECT  15.540 0.990 15.800 1.220 ;
        RECT  15.310 0.990 15.540 2.530 ;
        RECT  14.265 3.225 15.520 3.455 ;
        RECT  14.745 0.910 14.975 2.995 ;
        RECT  14.285 0.960 14.515 2.500 ;
        RECT  13.215 0.960 14.285 1.190 ;
        RECT  13.970 2.270 14.285 2.500 ;
        RECT  14.035 2.730 14.265 3.455 ;
        RECT  12.790 2.730 14.035 2.960 ;
        RECT  13.710 1.560 14.015 1.900 ;
        RECT  13.480 1.560 13.710 2.415 ;
        RECT  12.305 2.185 13.480 2.415 ;
        RECT  12.985 0.960 13.215 1.890 ;
        RECT  12.560 2.730 12.790 3.375 ;
        RECT  10.885 3.145 12.560 3.375 ;
        RECT  12.125 0.935 12.305 2.415 ;
        RECT  12.075 0.935 12.125 2.905 ;
        RECT  11.895 2.185 12.075 2.905 ;
        RECT  11.355 0.465 11.585 2.850 ;
        RECT  10.415 0.465 11.355 0.695 ;
        RECT  11.120 2.620 11.355 2.850 ;
        RECT  10.885 1.615 11.120 1.955 ;
        RECT  10.655 0.925 10.885 3.375 ;
        RECT  10.415 2.560 10.655 2.790 ;
        RECT  10.185 0.465 10.415 0.925 ;
        RECT  10.180 1.155 10.410 2.090 ;
        RECT  8.135 0.695 10.185 0.925 ;
        RECT  9.280 1.155 10.180 1.385 ;
        RECT  9.280 2.505 9.385 2.845 ;
        RECT  9.050 1.155 9.280 2.845 ;
        RECT  8.400 1.605 8.630 3.220 ;
        RECT  6.755 2.990 8.400 3.220 ;
        RECT  7.905 0.695 8.135 2.745 ;
        RECT  7.150 0.695 7.905 0.925 ;
        RECT  7.105 2.515 7.905 2.745 ;
        RECT  7.445 1.210 7.675 1.910 ;
        RECT  5.285 1.210 7.445 1.440 ;
        RECT  6.525 2.565 6.755 3.220 ;
        RECT  5.680 2.565 6.525 2.795 ;
        RECT  5.450 2.565 5.680 3.455 ;
        RECT  4.490 3.225 5.450 3.455 ;
        RECT  5.055 0.595 5.285 1.440 ;
        RECT  4.950 2.550 5.220 2.920 ;
        RECT  4.950 1.210 5.055 1.440 ;
        RECT  4.720 1.210 4.950 2.920 ;
        RECT  4.260 0.465 4.490 3.455 ;
        RECT  3.800 1.605 4.030 2.760 ;
        RECT  2.695 2.530 3.800 2.760 ;
        RECT  2.465 1.060 2.695 2.760 ;
        RECT  2.460 1.060 2.465 1.290 ;
        RECT  2.425 2.530 2.465 2.760 ;
        RECT  2.230 0.465 2.460 1.290 ;
        RECT  2.195 2.530 2.425 3.340 ;
        RECT  2.000 1.810 2.230 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFXD0BWP7T

MACRO SDFXD1BWP7T
    CLASS CORE ;
    FOREIGN SDFXD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 1.750 7.160 2.150 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.750 6.020 2.150 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.5040 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.060 1.075 18.340 2.560 ;
        RECT  17.925 1.075 18.060 1.305 ;
        RECT  17.640 2.330 18.060 2.560 ;
        RECT  17.695 0.480 17.925 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.130 0.470 19.460 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4248 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.735 3.360 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2241 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.760 9.940 2.710 ;
        RECT  9.510 1.760 9.660 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.700 -0.235 19.600 0.235 ;
        RECT  18.360 -0.235 18.700 0.810 ;
        RECT  15.570 -0.235 18.360 0.235 ;
        RECT  15.230 -0.235 15.570 0.465 ;
        RECT  13.550 -0.235 15.230 0.235 ;
        RECT  13.210 -0.235 13.550 0.730 ;
        RECT  9.955 -0.235 13.210 0.235 ;
        RECT  9.615 -0.235 9.955 0.465 ;
        RECT  8.835 -0.235 9.615 0.235 ;
        RECT  8.495 -0.235 8.835 0.465 ;
        RECT  6.115 -0.235 8.495 0.235 ;
        RECT  5.775 -0.235 6.115 0.840 ;
        RECT  3.795 -0.235 5.775 0.235 ;
        RECT  3.455 -0.235 3.795 1.145 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.700 3.685 19.600 4.155 ;
        RECT  18.360 3.250 18.700 4.155 ;
        RECT  16.560 3.685 18.360 4.155 ;
        RECT  16.220 3.250 16.560 4.155 ;
        RECT  13.560 3.685 16.220 4.155 ;
        RECT  13.200 3.190 13.560 4.155 ;
        RECT  10.000 3.685 13.200 4.155 ;
        RECT  9.660 3.455 10.000 4.155 ;
        RECT  8.865 3.685 9.660 4.155 ;
        RECT  8.525 3.455 8.865 4.155 ;
        RECT  6.140 3.685 8.525 4.155 ;
        RECT  5.910 3.025 6.140 4.155 ;
        RECT  3.825 3.685 5.910 4.155 ;
        RECT  3.485 3.020 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.655 1.600 18.885 3.020 ;
        RECT  17.410 2.790 18.655 3.020 ;
        RECT  16.030 0.465 17.460 0.695 ;
        RECT  17.225 1.020 17.410 3.020 ;
        RECT  17.180 1.020 17.225 3.380 ;
        RECT  16.490 1.020 17.180 1.250 ;
        RECT  16.995 2.565 17.180 3.380 ;
        RECT  16.720 1.565 16.950 2.310 ;
        RECT  16.490 2.080 16.720 2.310 ;
        RECT  16.260 1.020 16.490 1.830 ;
        RECT  16.260 2.080 16.490 2.995 ;
        RECT  15.775 1.600 16.260 1.830 ;
        RECT  14.975 2.765 16.260 2.995 ;
        RECT  15.800 0.465 16.030 1.220 ;
        RECT  15.540 2.300 15.810 2.530 ;
        RECT  15.540 0.990 15.800 1.220 ;
        RECT  15.310 0.990 15.540 2.530 ;
        RECT  14.265 3.225 15.520 3.455 ;
        RECT  14.745 0.910 14.975 2.995 ;
        RECT  14.285 0.960 14.515 2.500 ;
        RECT  13.215 0.960 14.285 1.190 ;
        RECT  13.970 2.270 14.285 2.500 ;
        RECT  14.035 2.730 14.265 3.455 ;
        RECT  12.790 2.730 14.035 2.960 ;
        RECT  13.710 1.560 14.015 1.900 ;
        RECT  13.480 1.560 13.710 2.415 ;
        RECT  12.305 2.185 13.480 2.415 ;
        RECT  12.985 0.960 13.215 1.890 ;
        RECT  12.560 2.730 12.790 3.375 ;
        RECT  10.885 3.145 12.560 3.375 ;
        RECT  12.125 0.935 12.305 2.415 ;
        RECT  12.075 0.935 12.125 2.905 ;
        RECT  11.895 2.185 12.075 2.905 ;
        RECT  11.355 0.465 11.585 2.850 ;
        RECT  10.415 0.465 11.355 0.695 ;
        RECT  11.120 2.620 11.355 2.850 ;
        RECT  10.885 1.615 11.120 1.955 ;
        RECT  10.655 0.925 10.885 3.375 ;
        RECT  10.415 2.560 10.655 2.790 ;
        RECT  10.185 0.465 10.415 0.925 ;
        RECT  10.180 1.155 10.410 2.090 ;
        RECT  8.135 0.695 10.185 0.925 ;
        RECT  9.280 1.155 10.180 1.385 ;
        RECT  9.280 2.505 9.385 2.845 ;
        RECT  9.050 1.155 9.280 2.845 ;
        RECT  8.400 1.605 8.630 3.220 ;
        RECT  6.755 2.990 8.400 3.220 ;
        RECT  7.905 0.695 8.135 2.745 ;
        RECT  7.150 0.695 7.905 0.925 ;
        RECT  7.105 2.515 7.905 2.745 ;
        RECT  7.445 1.210 7.675 1.910 ;
        RECT  5.285 1.210 7.445 1.440 ;
        RECT  6.525 2.565 6.755 3.220 ;
        RECT  5.680 2.565 6.525 2.795 ;
        RECT  5.450 2.565 5.680 3.455 ;
        RECT  4.490 3.225 5.450 3.455 ;
        RECT  5.055 0.595 5.285 1.440 ;
        RECT  4.950 2.550 5.220 2.920 ;
        RECT  4.950 1.210 5.055 1.440 ;
        RECT  4.720 1.210 4.950 2.920 ;
        RECT  4.260 0.465 4.490 3.455 ;
        RECT  3.800 1.605 4.030 2.760 ;
        RECT  2.695 2.530 3.800 2.760 ;
        RECT  2.465 1.060 2.695 2.760 ;
        RECT  2.460 1.060 2.465 1.290 ;
        RECT  2.425 2.530 2.465 2.760 ;
        RECT  2.230 0.465 2.460 1.290 ;
        RECT  2.195 2.530 2.425 3.340 ;
        RECT  2.000 1.810 2.230 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFXD1BWP7T

MACRO SDFXD2BWP7T
    CLASS CORE ;
    FOREIGN SDFXD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 1.750 7.160 2.150 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.750 6.020 2.150 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.5040 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SA
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.600 0.465 18.945 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.325 1.055 20.580 2.690 ;
        RECT  20.300 0.465 20.325 3.310 ;
        RECT  20.090 0.465 20.300 1.285 ;
        RECT  20.095 2.460 20.300 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4248 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.735 3.360 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2241 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.760 9.940 2.710 ;
        RECT  9.510 1.760 9.660 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.045 -0.235 21.280 0.235 ;
        RECT  20.815 -0.235 21.045 1.245 ;
        RECT  19.660 -0.235 20.815 0.235 ;
        RECT  19.320 -0.235 19.660 1.180 ;
        RECT  18.180 -0.235 19.320 0.235 ;
        RECT  17.840 -0.235 18.180 0.465 ;
        RECT  16.565 -0.235 17.840 0.235 ;
        RECT  16.225 -0.235 16.565 0.465 ;
        RECT  13.550 -0.235 16.225 0.235 ;
        RECT  13.210 -0.235 13.550 0.730 ;
        RECT  9.955 -0.235 13.210 0.235 ;
        RECT  9.615 -0.235 9.955 0.465 ;
        RECT  8.835 -0.235 9.615 0.235 ;
        RECT  8.495 -0.235 8.835 0.465 ;
        RECT  6.115 -0.235 8.495 0.235 ;
        RECT  5.775 -0.235 6.115 0.840 ;
        RECT  3.795 -0.235 5.775 0.235 ;
        RECT  3.455 -0.235 3.795 1.145 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.045 3.685 21.280 4.155 ;
        RECT  20.815 2.255 21.045 4.155 ;
        RECT  19.660 3.685 20.815 4.155 ;
        RECT  19.320 3.250 19.660 4.155 ;
        RECT  18.145 3.685 19.320 4.155 ;
        RECT  17.805 3.250 18.145 4.155 ;
        RECT  16.615 3.685 17.805 4.155 ;
        RECT  16.275 3.250 16.615 4.155 ;
        RECT  13.560 3.685 16.275 4.155 ;
        RECT  13.200 3.190 13.560 4.155 ;
        RECT  10.000 3.685 13.200 4.155 ;
        RECT  9.660 3.455 10.000 4.155 ;
        RECT  8.865 3.685 9.660 4.155 ;
        RECT  8.525 3.455 8.865 4.155 ;
        RECT  6.140 3.685 8.525 4.155 ;
        RECT  5.910 3.025 6.140 4.155 ;
        RECT  3.825 3.685 5.910 4.155 ;
        RECT  3.485 3.020 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.615 1.600 19.845 3.010 ;
        RECT  17.595 2.780 19.615 3.010 ;
        RECT  18.130 0.695 18.360 1.940 ;
        RECT  16.030 0.695 18.130 0.925 ;
        RECT  17.365 1.155 17.595 3.010 ;
        RECT  16.545 1.155 17.365 1.385 ;
        RECT  17.325 2.565 17.365 3.010 ;
        RECT  17.095 2.565 17.325 3.380 ;
        RECT  16.840 1.675 17.070 2.310 ;
        RECT  16.570 2.080 16.840 2.310 ;
        RECT  16.340 2.080 16.570 2.995 ;
        RECT  16.315 1.155 16.545 1.830 ;
        RECT  14.975 2.765 16.340 2.995 ;
        RECT  15.765 1.600 16.315 1.830 ;
        RECT  15.800 0.695 16.030 1.220 ;
        RECT  15.500 2.300 15.810 2.530 ;
        RECT  15.500 0.990 15.800 1.220 ;
        RECT  15.270 0.990 15.500 2.530 ;
        RECT  14.265 3.225 15.465 3.455 ;
        RECT  14.745 0.910 14.975 2.995 ;
        RECT  14.285 0.960 14.515 2.500 ;
        RECT  13.215 0.960 14.285 1.190 ;
        RECT  13.970 2.270 14.285 2.500 ;
        RECT  14.035 2.730 14.265 3.455 ;
        RECT  12.790 2.730 14.035 2.960 ;
        RECT  13.710 1.560 14.015 1.900 ;
        RECT  13.480 1.560 13.710 2.415 ;
        RECT  12.305 2.185 13.480 2.415 ;
        RECT  12.985 0.960 13.215 1.890 ;
        RECT  12.560 2.730 12.790 3.375 ;
        RECT  10.885 3.145 12.560 3.375 ;
        RECT  12.125 0.935 12.305 2.415 ;
        RECT  12.075 0.935 12.125 2.905 ;
        RECT  11.895 2.185 12.075 2.905 ;
        RECT  11.355 0.465 11.585 2.850 ;
        RECT  10.415 0.465 11.355 0.695 ;
        RECT  11.120 2.620 11.355 2.850 ;
        RECT  10.885 1.615 11.120 1.955 ;
        RECT  10.655 0.925 10.885 3.375 ;
        RECT  10.415 2.560 10.655 2.790 ;
        RECT  10.185 0.465 10.415 0.925 ;
        RECT  10.180 1.155 10.410 2.090 ;
        RECT  8.135 0.695 10.185 0.925 ;
        RECT  9.280 1.155 10.180 1.385 ;
        RECT  9.280 2.505 9.385 2.845 ;
        RECT  9.050 1.155 9.280 2.845 ;
        RECT  8.400 1.605 8.630 3.220 ;
        RECT  6.755 2.990 8.400 3.220 ;
        RECT  7.905 0.695 8.135 2.745 ;
        RECT  7.150 0.695 7.905 0.925 ;
        RECT  7.105 2.515 7.905 2.745 ;
        RECT  7.445 1.210 7.675 1.910 ;
        RECT  5.285 1.210 7.445 1.440 ;
        RECT  6.525 2.565 6.755 3.220 ;
        RECT  5.680 2.565 6.525 2.795 ;
        RECT  5.450 2.565 5.680 3.455 ;
        RECT  4.490 3.225 5.450 3.455 ;
        RECT  5.055 0.595 5.285 1.440 ;
        RECT  4.950 2.550 5.220 2.920 ;
        RECT  4.950 1.210 5.055 1.440 ;
        RECT  4.720 1.210 4.950 2.920 ;
        RECT  4.260 0.465 4.490 3.455 ;
        RECT  3.800 1.605 4.030 2.760 ;
        RECT  2.695 2.530 3.800 2.760 ;
        RECT  2.465 1.060 2.695 2.760 ;
        RECT  2.460 1.060 2.465 1.290 ;
        RECT  2.425 2.530 2.465 2.760 ;
        RECT  2.230 0.465 2.460 1.290 ;
        RECT  2.195 2.530 2.425 3.340 ;
        RECT  2.000 1.810 2.230 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFXD2BWP7T

MACRO SDFXQD0BWP7T
    CLASS CORE ;
    FOREIGN SDFXQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 1.750 7.160 2.150 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.750 6.020 2.150 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.5040 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 0.5925 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.570 0.510 18.900 3.405 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4248 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.735 3.360 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2241 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.760 9.940 2.710 ;
        RECT  9.510 1.760 9.660 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.045 -0.235 19.040 0.235 ;
        RECT  17.815 -0.235 18.045 0.860 ;
        RECT  16.665 -0.235 17.815 0.235 ;
        RECT  16.325 -0.235 16.665 0.740 ;
        RECT  13.550 -0.235 16.325 0.235 ;
        RECT  13.210 -0.235 13.550 0.730 ;
        RECT  9.955 -0.235 13.210 0.235 ;
        RECT  9.615 -0.235 9.955 0.465 ;
        RECT  8.835 -0.235 9.615 0.235 ;
        RECT  8.495 -0.235 8.835 0.465 ;
        RECT  6.115 -0.235 8.495 0.235 ;
        RECT  5.775 -0.235 6.115 0.840 ;
        RECT  3.795 -0.235 5.775 0.235 ;
        RECT  3.455 -0.235 3.795 1.145 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.045 3.685 19.040 4.155 ;
        RECT  17.815 3.065 18.045 4.155 ;
        RECT  16.675 3.685 17.815 4.155 ;
        RECT  16.335 3.250 16.675 4.155 ;
        RECT  13.560 3.685 16.335 4.155 ;
        RECT  13.200 3.190 13.560 4.155 ;
        RECT  10.000 3.685 13.200 4.155 ;
        RECT  9.660 3.455 10.000 4.155 ;
        RECT  8.865 3.685 9.660 4.155 ;
        RECT  8.525 3.455 8.865 4.155 ;
        RECT  6.140 3.685 8.525 4.155 ;
        RECT  5.910 3.025 6.140 4.155 ;
        RECT  3.825 3.685 5.910 4.155 ;
        RECT  3.485 3.020 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.585 1.670 18.305 2.010 ;
        RECT  17.355 1.040 17.585 2.795 ;
        RECT  17.340 1.040 17.355 1.270 ;
        RECT  17.340 2.565 17.355 2.795 ;
        RECT  17.110 0.495 17.340 1.270 ;
        RECT  17.110 2.565 17.340 3.380 ;
        RECT  16.885 1.565 17.115 2.310 ;
        RECT  16.505 1.040 17.110 1.270 ;
        RECT  16.605 2.080 16.885 2.310 ;
        RECT  16.375 2.080 16.605 2.995 ;
        RECT  16.275 1.040 16.505 1.830 ;
        RECT  15.015 2.765 16.375 2.995 ;
        RECT  15.890 1.600 16.275 1.830 ;
        RECT  15.575 2.300 15.870 2.530 ;
        RECT  15.575 0.990 15.830 1.220 ;
        RECT  14.265 3.225 15.580 3.455 ;
        RECT  15.345 0.990 15.575 2.530 ;
        RECT  14.785 0.910 15.015 2.995 ;
        RECT  14.285 0.960 14.515 2.500 ;
        RECT  13.215 0.960 14.285 1.190 ;
        RECT  13.970 2.270 14.285 2.500 ;
        RECT  14.035 2.730 14.265 3.455 ;
        RECT  12.790 2.730 14.035 2.960 ;
        RECT  13.710 1.560 14.015 1.900 ;
        RECT  13.480 1.560 13.710 2.415 ;
        RECT  12.305 2.185 13.480 2.415 ;
        RECT  12.985 0.960 13.215 1.890 ;
        RECT  12.560 2.730 12.790 3.375 ;
        RECT  10.885 3.145 12.560 3.375 ;
        RECT  12.125 0.935 12.305 2.415 ;
        RECT  12.075 0.935 12.125 2.905 ;
        RECT  11.895 2.185 12.075 2.905 ;
        RECT  11.355 0.465 11.585 2.850 ;
        RECT  10.415 0.465 11.355 0.695 ;
        RECT  11.120 2.620 11.355 2.850 ;
        RECT  10.885 1.615 11.120 1.955 ;
        RECT  10.655 0.925 10.885 3.375 ;
        RECT  10.415 2.560 10.655 2.790 ;
        RECT  10.185 0.465 10.415 0.925 ;
        RECT  10.180 1.155 10.410 2.090 ;
        RECT  8.135 0.695 10.185 0.925 ;
        RECT  9.280 1.155 10.180 1.385 ;
        RECT  9.280 2.505 9.385 2.845 ;
        RECT  9.050 1.155 9.280 2.845 ;
        RECT  8.400 1.605 8.630 3.220 ;
        RECT  6.755 2.990 8.400 3.220 ;
        RECT  7.905 0.695 8.135 2.745 ;
        RECT  7.150 0.695 7.905 0.925 ;
        RECT  7.105 2.515 7.905 2.745 ;
        RECT  7.445 1.210 7.675 1.910 ;
        RECT  5.285 1.210 7.445 1.440 ;
        RECT  6.525 2.565 6.755 3.220 ;
        RECT  5.680 2.565 6.525 2.795 ;
        RECT  5.450 2.565 5.680 3.455 ;
        RECT  4.490 3.225 5.450 3.455 ;
        RECT  5.055 0.595 5.285 1.440 ;
        RECT  4.950 2.550 5.220 2.920 ;
        RECT  4.950 1.210 5.055 1.440 ;
        RECT  4.720 1.210 4.950 2.920 ;
        RECT  4.260 0.465 4.490 3.455 ;
        RECT  3.800 1.605 4.030 2.760 ;
        RECT  2.695 2.530 3.800 2.760 ;
        RECT  2.465 1.060 2.695 2.760 ;
        RECT  2.460 1.060 2.465 1.290 ;
        RECT  2.425 2.530 2.465 2.760 ;
        RECT  2.230 0.465 2.460 1.290 ;
        RECT  2.195 2.530 2.425 3.340 ;
        RECT  2.000 1.810 2.230 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFXQD0BWP7T

MACRO SDFXQD1BWP7T
    CLASS CORE ;
    FOREIGN SDFXQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 1.750 7.160 2.150 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.750 6.020 2.150 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.5040 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 1.1850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.570 0.470 18.900 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4248 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.735 3.360 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2241 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.760 9.940 2.710 ;
        RECT  9.510 1.760 9.660 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.045 -0.235 19.040 0.235 ;
        RECT  17.815 -0.235 18.045 1.255 ;
        RECT  16.665 -0.235 17.815 0.235 ;
        RECT  16.325 -0.235 16.665 0.670 ;
        RECT  13.550 -0.235 16.325 0.235 ;
        RECT  13.210 -0.235 13.550 0.730 ;
        RECT  9.955 -0.235 13.210 0.235 ;
        RECT  9.615 -0.235 9.955 0.465 ;
        RECT  8.835 -0.235 9.615 0.235 ;
        RECT  8.495 -0.235 8.835 0.465 ;
        RECT  6.115 -0.235 8.495 0.235 ;
        RECT  5.775 -0.235 6.115 0.840 ;
        RECT  3.795 -0.235 5.775 0.235 ;
        RECT  3.455 -0.235 3.795 1.145 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.045 3.685 19.040 4.155 ;
        RECT  17.815 2.255 18.045 4.155 ;
        RECT  16.675 3.685 17.815 4.155 ;
        RECT  16.335 3.250 16.675 4.155 ;
        RECT  13.560 3.685 16.335 4.155 ;
        RECT  13.200 3.190 13.560 4.155 ;
        RECT  10.000 3.685 13.200 4.155 ;
        RECT  9.660 3.455 10.000 4.155 ;
        RECT  8.865 3.685 9.660 4.155 ;
        RECT  8.525 3.455 8.865 4.155 ;
        RECT  6.140 3.685 8.525 4.155 ;
        RECT  5.910 3.025 6.140 4.155 ;
        RECT  3.825 3.685 5.910 4.155 ;
        RECT  3.485 3.020 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.585 1.600 18.305 1.940 ;
        RECT  17.355 1.020 17.585 2.795 ;
        RECT  17.340 1.020 17.355 1.250 ;
        RECT  17.340 2.565 17.355 2.795 ;
        RECT  17.110 0.495 17.340 1.250 ;
        RECT  17.110 2.565 17.340 3.380 ;
        RECT  16.885 1.565 17.115 2.310 ;
        RECT  16.505 1.020 17.110 1.250 ;
        RECT  16.605 2.080 16.885 2.310 ;
        RECT  16.375 2.080 16.605 2.995 ;
        RECT  16.275 1.020 16.505 1.830 ;
        RECT  15.015 2.765 16.375 2.995 ;
        RECT  15.890 1.600 16.275 1.830 ;
        RECT  15.575 2.300 15.870 2.530 ;
        RECT  15.575 0.990 15.830 1.220 ;
        RECT  14.265 3.225 15.580 3.455 ;
        RECT  15.345 0.990 15.575 2.530 ;
        RECT  14.785 0.910 15.015 2.995 ;
        RECT  14.285 0.960 14.515 2.500 ;
        RECT  13.215 0.960 14.285 1.190 ;
        RECT  13.970 2.270 14.285 2.500 ;
        RECT  14.035 2.730 14.265 3.455 ;
        RECT  12.790 2.730 14.035 2.960 ;
        RECT  13.710 1.560 14.015 1.900 ;
        RECT  13.480 1.560 13.710 2.415 ;
        RECT  12.305 2.185 13.480 2.415 ;
        RECT  12.985 0.960 13.215 1.890 ;
        RECT  12.560 2.730 12.790 3.375 ;
        RECT  10.885 3.145 12.560 3.375 ;
        RECT  12.125 0.935 12.305 2.415 ;
        RECT  12.075 0.935 12.125 2.905 ;
        RECT  11.895 2.185 12.075 2.905 ;
        RECT  11.355 0.465 11.585 2.850 ;
        RECT  10.415 0.465 11.355 0.695 ;
        RECT  11.120 2.620 11.355 2.850 ;
        RECT  10.885 1.615 11.120 1.955 ;
        RECT  10.655 0.925 10.885 3.375 ;
        RECT  10.415 2.560 10.655 2.790 ;
        RECT  10.185 0.465 10.415 0.925 ;
        RECT  10.180 1.155 10.410 2.090 ;
        RECT  8.135 0.695 10.185 0.925 ;
        RECT  9.280 1.155 10.180 1.385 ;
        RECT  9.280 2.505 9.385 2.845 ;
        RECT  9.050 1.155 9.280 2.845 ;
        RECT  8.400 1.605 8.630 3.220 ;
        RECT  6.755 2.990 8.400 3.220 ;
        RECT  7.905 0.695 8.135 2.745 ;
        RECT  7.150 0.695 7.905 0.925 ;
        RECT  7.105 2.515 7.905 2.745 ;
        RECT  7.445 1.210 7.675 1.910 ;
        RECT  5.285 1.210 7.445 1.440 ;
        RECT  6.525 2.565 6.755 3.220 ;
        RECT  5.680 2.565 6.525 2.795 ;
        RECT  5.450 2.565 5.680 3.455 ;
        RECT  4.490 3.225 5.450 3.455 ;
        RECT  5.055 0.595 5.285 1.440 ;
        RECT  4.950 2.550 5.220 2.920 ;
        RECT  4.950 1.210 5.055 1.440 ;
        RECT  4.720 1.210 4.950 2.920 ;
        RECT  4.260 0.465 4.490 3.455 ;
        RECT  3.800 1.605 4.030 2.760 ;
        RECT  2.695 2.530 3.800 2.760 ;
        RECT  2.465 1.060 2.695 2.760 ;
        RECT  2.460 1.060 2.465 1.290 ;
        RECT  2.425 2.530 2.465 2.760 ;
        RECT  2.230 0.465 2.460 1.290 ;
        RECT  2.195 2.530 2.425 3.340 ;
        RECT  2.000 1.810 2.230 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFXQD1BWP7T

MACRO SDFXQD2BWP7T
    CLASS CORE ;
    FOREIGN SDFXQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 1.750 7.160 2.150 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4860 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 1.750 6.020 2.150 ;
        END
    END SE
    PIN SA
        ANTENNAGATEAREA 0.5040 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 1.590 0.980 2.710 ;
        END
    END SA
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.645 1.045 18.900 2.730 ;
        RECT  18.620 0.465 18.645 3.310 ;
        RECT  18.415 0.465 18.620 1.280 ;
        RECT  18.415 2.500 18.620 3.310 ;
        END
    END Q
    PIN DB
        ANTENNAGATEAREA 0.4248 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.735 3.360 2.150 ;
        RECT  2.940 1.210 3.220 2.150 ;
        END
    END DB
    PIN DA
        ANTENNAGATEAREA 0.2241 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.590 1.540 2.710 ;
        END
    END DA
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.760 9.940 2.710 ;
        RECT  9.510 1.760 9.660 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.365 -0.235 19.600 0.235 ;
        RECT  19.135 -0.235 19.365 1.230 ;
        RECT  17.925 -0.235 19.135 0.235 ;
        RECT  17.695 -0.235 17.925 1.255 ;
        RECT  16.470 -0.235 17.695 0.235 ;
        RECT  16.130 -0.235 16.470 0.745 ;
        RECT  13.550 -0.235 16.130 0.235 ;
        RECT  13.210 -0.235 13.550 0.730 ;
        RECT  9.955 -0.235 13.210 0.235 ;
        RECT  9.615 -0.235 9.955 0.465 ;
        RECT  8.835 -0.235 9.615 0.235 ;
        RECT  8.495 -0.235 8.835 0.465 ;
        RECT  6.115 -0.235 8.495 0.235 ;
        RECT  5.775 -0.235 6.115 0.840 ;
        RECT  3.795 -0.235 5.775 0.235 ;
        RECT  3.455 -0.235 3.795 1.145 ;
        RECT  1.240 -0.235 3.455 0.235 ;
        RECT  0.900 -0.235 1.240 0.840 ;
        RECT  0.000 -0.235 0.900 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.365 3.685 19.600 4.155 ;
        RECT  19.135 2.255 19.365 4.155 ;
        RECT  17.925 3.685 19.135 4.155 ;
        RECT  17.695 2.255 17.925 4.155 ;
        RECT  16.490 3.685 17.695 4.155 ;
        RECT  16.150 2.545 16.490 4.155 ;
        RECT  13.560 3.685 16.150 4.155 ;
        RECT  13.200 3.190 13.560 4.155 ;
        RECT  10.000 3.685 13.200 4.155 ;
        RECT  9.660 3.455 10.000 4.155 ;
        RECT  8.865 3.685 9.660 4.155 ;
        RECT  8.525 3.455 8.865 4.155 ;
        RECT  6.140 3.685 8.525 4.155 ;
        RECT  5.910 3.025 6.140 4.155 ;
        RECT  3.825 3.685 5.910 4.155 ;
        RECT  3.485 3.020 3.825 4.155 ;
        RECT  1.240 3.685 3.485 4.155 ;
        RECT  0.900 2.945 1.240 4.155 ;
        RECT  0.000 3.685 0.900 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.460 1.600 18.305 1.940 ;
        RECT  17.230 1.020 17.460 2.795 ;
        RECT  17.205 1.020 17.230 1.250 ;
        RECT  17.205 2.565 17.230 2.795 ;
        RECT  16.975 0.495 17.205 1.250 ;
        RECT  16.975 2.565 17.205 3.380 ;
        RECT  16.750 1.590 16.980 2.310 ;
        RECT  16.320 1.020 16.975 1.250 ;
        RECT  15.015 2.080 16.750 2.310 ;
        RECT  16.090 1.020 16.320 1.830 ;
        RECT  15.715 1.600 16.090 1.830 ;
        RECT  14.265 3.225 15.465 3.455 ;
        RECT  14.785 0.910 15.015 2.850 ;
        RECT  14.285 0.960 14.515 2.500 ;
        RECT  13.215 0.960 14.285 1.190 ;
        RECT  13.970 2.270 14.285 2.500 ;
        RECT  14.035 2.730 14.265 3.455 ;
        RECT  12.790 2.730 14.035 2.960 ;
        RECT  13.710 1.560 14.015 1.900 ;
        RECT  13.480 1.560 13.710 2.415 ;
        RECT  12.305 2.185 13.480 2.415 ;
        RECT  12.985 0.960 13.215 1.890 ;
        RECT  12.560 2.730 12.790 3.375 ;
        RECT  10.885 3.145 12.560 3.375 ;
        RECT  12.125 0.935 12.305 2.415 ;
        RECT  12.075 0.935 12.125 2.905 ;
        RECT  11.895 2.185 12.075 2.905 ;
        RECT  11.355 0.465 11.585 2.850 ;
        RECT  10.415 0.465 11.355 0.695 ;
        RECT  11.120 2.620 11.355 2.850 ;
        RECT  10.885 1.615 11.120 1.955 ;
        RECT  10.655 0.925 10.885 3.375 ;
        RECT  10.415 2.560 10.655 2.790 ;
        RECT  10.185 0.465 10.415 0.925 ;
        RECT  10.180 1.155 10.410 2.090 ;
        RECT  8.135 0.695 10.185 0.925 ;
        RECT  9.280 1.155 10.180 1.385 ;
        RECT  9.280 2.505 9.385 2.845 ;
        RECT  9.050 1.155 9.280 2.845 ;
        RECT  8.400 1.605 8.630 3.220 ;
        RECT  6.755 2.990 8.400 3.220 ;
        RECT  7.905 0.695 8.135 2.745 ;
        RECT  7.150 0.695 7.905 0.925 ;
        RECT  7.105 2.515 7.905 2.745 ;
        RECT  7.445 1.210 7.675 1.910 ;
        RECT  5.285 1.210 7.445 1.440 ;
        RECT  6.525 2.565 6.755 3.220 ;
        RECT  5.680 2.565 6.525 2.795 ;
        RECT  5.450 2.565 5.680 3.455 ;
        RECT  4.490 3.225 5.450 3.455 ;
        RECT  5.055 0.595 5.285 1.440 ;
        RECT  4.950 2.550 5.220 2.920 ;
        RECT  4.950 1.210 5.055 1.440 ;
        RECT  4.720 1.210 4.950 2.920 ;
        RECT  4.260 0.465 4.490 3.455 ;
        RECT  3.800 1.605 4.030 2.760 ;
        RECT  2.695 2.530 3.800 2.760 ;
        RECT  2.465 1.060 2.695 2.760 ;
        RECT  2.460 1.060 2.465 1.290 ;
        RECT  2.425 2.530 2.465 2.760 ;
        RECT  2.230 0.465 2.460 1.290 ;
        RECT  2.195 2.530 2.425 3.340 ;
        RECT  2.000 1.810 2.230 2.150 ;
        RECT  1.770 1.130 2.000 2.150 ;
        RECT  0.465 1.130 1.770 1.360 ;
        RECT  0.345 2.950 0.520 3.180 ;
        RECT  0.345 0.595 0.465 1.360 ;
        RECT  0.235 0.595 0.345 3.180 ;
        RECT  0.115 1.130 0.235 3.180 ;
    END
END SDFXQD2BWP7T

MACRO SEDFCND0BWP7T
    CLASS CORE ;
    FOREIGN SEDFCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.180 1.075 19.460 2.560 ;
        RECT  19.045 1.075 19.180 1.305 ;
        RECT  18.760 2.330 19.180 2.560 ;
        RECT  18.815 0.505 19.045 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.250 0.505 20.580 2.715 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.820 8.340 2.115 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.3942 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.160 2.395 17.275 2.625 ;
        RECT  16.930 2.395 17.160 3.455 ;
        RECT  14.950 3.225 16.930 3.455 ;
        RECT  14.720 2.730 14.950 3.455 ;
        RECT  13.790 2.730 14.720 2.960 ;
        RECT  13.560 2.730 13.790 3.270 ;
        RECT  11.785 2.940 13.560 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.820 -0.235 20.720 0.235 ;
        RECT  19.480 -0.235 19.820 0.790 ;
        RECT  16.090 -0.235 19.480 0.235 ;
        RECT  15.750 -0.235 16.090 0.465 ;
        RECT  12.815 -0.235 15.750 0.235 ;
        RECT  12.475 -0.235 12.815 0.730 ;
        RECT  8.670 -0.235 12.475 0.235 ;
        RECT  8.330 -0.235 8.670 0.465 ;
        RECT  4.035 -0.235 8.330 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.780 3.685 20.720 4.155 ;
        RECT  19.440 3.355 19.780 4.155 ;
        RECT  18.560 3.685 19.440 4.155 ;
        RECT  18.220 3.455 18.560 4.155 ;
        RECT  14.480 3.685 18.220 4.155 ;
        RECT  14.140 3.190 14.480 4.155 ;
        RECT  8.205 3.685 14.140 4.155 ;
        RECT  7.865 3.440 8.205 4.155 ;
        RECT  3.995 3.685 7.865 4.155 ;
        RECT  3.635 2.950 3.995 4.155 ;
        RECT  1.290 3.685 3.635 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.775 1.600 20.005 3.020 ;
        RECT  18.495 2.790 19.775 3.020 ;
        RECT  16.770 0.465 18.580 0.695 ;
        RECT  18.265 1.020 18.495 3.020 ;
        RECT  17.410 1.020 18.265 1.250 ;
        RECT  17.740 2.390 18.265 2.620 ;
        RECT  17.755 1.565 17.985 2.160 ;
        RECT  16.700 1.930 17.755 2.160 ;
        RECT  17.510 2.390 17.740 3.200 ;
        RECT  17.180 1.020 17.410 1.700 ;
        RECT  16.200 1.470 17.180 1.700 ;
        RECT  16.540 0.465 16.770 1.180 ;
        RECT  16.470 1.930 16.700 2.995 ;
        RECT  15.920 0.950 16.540 1.180 ;
        RECT  15.415 2.765 16.470 2.995 ;
        RECT  15.920 2.305 16.190 2.535 ;
        RECT  15.690 0.950 15.920 2.535 ;
        RECT  15.165 0.950 15.690 1.220 ;
        RECT  15.185 1.615 15.415 2.995 ;
        RECT  14.610 1.615 15.185 1.845 ;
        RECT  14.935 0.465 15.165 1.220 ;
        RECT  13.275 0.465 14.935 0.695 ;
        RECT  14.380 0.990 14.610 1.845 ;
        RECT  13.990 2.270 14.505 2.500 ;
        RECT  14.150 0.990 14.380 1.220 ;
        RECT  13.760 1.420 13.990 2.500 ;
        RECT  13.735 1.420 13.760 1.650 ;
        RECT  13.505 0.925 13.735 1.650 ;
        RECT  12.725 1.420 13.505 1.650 ;
        RECT  13.055 1.880 13.395 2.200 ;
        RECT  13.045 0.465 13.275 1.190 ;
        RECT  11.545 2.440 13.205 2.670 ;
        RECT  11.025 1.970 13.055 2.200 ;
        RECT  11.780 0.960 13.045 1.190 ;
        RECT  12.385 1.420 12.725 1.740 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  9.135 0.465 11.550 0.695 ;
        RECT  11.020 1.970 11.025 2.725 ;
        RECT  10.790 0.935 11.020 2.725 ;
        RECT  10.255 0.990 10.390 2.865 ;
        RECT  10.155 0.990 10.255 3.210 ;
        RECT  9.965 0.990 10.155 1.220 ;
        RECT  10.025 2.525 10.155 3.210 ;
        RECT  7.775 2.980 10.025 3.210 ;
        RECT  9.725 1.805 9.925 2.035 ;
        RECT  9.495 1.115 9.725 2.670 ;
        RECT  9.265 1.115 9.495 1.345 ;
        RECT  9.270 2.440 9.495 2.670 ;
        RECT  9.005 1.800 9.200 2.040 ;
        RECT  8.905 0.465 9.135 0.925 ;
        RECT  8.775 1.155 9.005 2.725 ;
        RECT  7.700 0.695 8.905 0.925 ;
        RECT  7.940 1.155 8.775 1.385 ;
        RECT  8.005 2.380 8.775 2.725 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.470 0.695 7.700 1.590 ;
        RECT  6.215 2.555 7.545 2.785 ;
        RECT  6.935 1.360 7.470 1.590 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.890 0.505 7.230 1.130 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  6.705 1.360 6.935 2.220 ;
        RECT  4.540 0.505 6.890 0.735 ;
        RECT  5.985 0.965 6.215 2.785 ;
        RECT  4.585 0.965 5.985 1.195 ;
        RECT  5.725 2.555 5.985 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.415 0.965 4.585 1.250 ;
        RECT  3.575 1.020 4.415 1.250 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.590 0.465 2.960 ;
    END
END SEDFCND0BWP7T

MACRO SEDFCND1BWP7T
    CLASS CORE ;
    FOREIGN SEDFCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.9672 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.180 1.075 19.460 2.560 ;
        RECT  19.045 1.075 19.180 1.305 ;
        RECT  18.760 2.330 19.180 2.560 ;
        RECT  18.815 0.480 19.045 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.250 0.470 20.580 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.820 8.340 2.115 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.3942 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.160 2.395 17.275 2.625 ;
        RECT  16.930 2.395 17.160 3.455 ;
        RECT  14.950 3.225 16.930 3.455 ;
        RECT  14.720 2.730 14.950 3.455 ;
        RECT  13.790 2.730 14.720 2.960 ;
        RECT  13.560 2.730 13.790 3.270 ;
        RECT  11.785 2.940 13.560 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.820 -0.235 20.720 0.235 ;
        RECT  19.480 -0.235 19.820 0.810 ;
        RECT  16.090 -0.235 19.480 0.235 ;
        RECT  15.750 -0.235 16.090 0.465 ;
        RECT  12.815 -0.235 15.750 0.235 ;
        RECT  12.475 -0.235 12.815 0.730 ;
        RECT  8.670 -0.235 12.475 0.235 ;
        RECT  8.330 -0.235 8.670 0.465 ;
        RECT  4.035 -0.235 8.330 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.820 3.685 20.720 4.155 ;
        RECT  19.480 3.250 19.820 4.155 ;
        RECT  18.560 3.685 19.480 4.155 ;
        RECT  18.220 3.455 18.560 4.155 ;
        RECT  14.480 3.685 18.220 4.155 ;
        RECT  14.140 3.190 14.480 4.155 ;
        RECT  8.205 3.685 14.140 4.155 ;
        RECT  7.865 3.440 8.205 4.155 ;
        RECT  3.995 3.685 7.865 4.155 ;
        RECT  3.635 2.950 3.995 4.155 ;
        RECT  1.290 3.685 3.635 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.775 1.600 20.005 3.020 ;
        RECT  18.495 2.790 19.775 3.020 ;
        RECT  16.770 0.465 18.580 0.695 ;
        RECT  18.265 1.020 18.495 3.020 ;
        RECT  17.410 1.020 18.265 1.250 ;
        RECT  17.740 2.390 18.265 2.620 ;
        RECT  17.755 1.565 17.985 2.160 ;
        RECT  16.700 1.930 17.755 2.160 ;
        RECT  17.510 2.390 17.740 3.200 ;
        RECT  17.180 1.020 17.410 1.700 ;
        RECT  16.200 1.470 17.180 1.700 ;
        RECT  16.540 0.465 16.770 1.180 ;
        RECT  16.470 1.930 16.700 2.995 ;
        RECT  15.920 0.950 16.540 1.180 ;
        RECT  15.415 2.765 16.470 2.995 ;
        RECT  15.920 2.305 16.190 2.535 ;
        RECT  15.690 0.950 15.920 2.535 ;
        RECT  15.165 0.950 15.690 1.220 ;
        RECT  15.185 1.615 15.415 2.995 ;
        RECT  14.610 1.615 15.185 1.845 ;
        RECT  14.935 0.465 15.165 1.220 ;
        RECT  13.275 0.465 14.935 0.695 ;
        RECT  14.380 0.990 14.610 1.845 ;
        RECT  13.990 2.270 14.505 2.500 ;
        RECT  14.150 0.990 14.380 1.220 ;
        RECT  13.760 1.420 13.990 2.500 ;
        RECT  13.735 1.420 13.760 1.650 ;
        RECT  13.505 0.925 13.735 1.650 ;
        RECT  12.725 1.420 13.505 1.650 ;
        RECT  13.055 1.880 13.395 2.200 ;
        RECT  13.045 0.465 13.275 1.190 ;
        RECT  11.545 2.440 13.205 2.670 ;
        RECT  11.025 1.970 13.055 2.200 ;
        RECT  11.780 0.960 13.045 1.190 ;
        RECT  12.385 1.420 12.725 1.740 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  9.135 0.465 11.550 0.695 ;
        RECT  11.020 1.970 11.025 2.725 ;
        RECT  10.790 0.935 11.020 2.725 ;
        RECT  10.255 0.990 10.390 2.865 ;
        RECT  10.155 0.990 10.255 3.210 ;
        RECT  9.965 0.990 10.155 1.220 ;
        RECT  10.025 2.525 10.155 3.210 ;
        RECT  7.775 2.980 10.025 3.210 ;
        RECT  9.725 1.805 9.925 2.035 ;
        RECT  9.495 1.115 9.725 2.670 ;
        RECT  9.265 1.115 9.495 1.345 ;
        RECT  9.270 2.440 9.495 2.670 ;
        RECT  9.005 1.800 9.200 2.040 ;
        RECT  8.905 0.465 9.135 0.925 ;
        RECT  8.775 1.155 9.005 2.725 ;
        RECT  7.700 0.695 8.905 0.925 ;
        RECT  7.940 1.155 8.775 1.385 ;
        RECT  8.005 2.380 8.775 2.725 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.470 0.695 7.700 1.590 ;
        RECT  6.215 2.555 7.545 2.785 ;
        RECT  6.935 1.360 7.470 1.590 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.890 0.505 7.230 1.130 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  6.705 1.360 6.935 2.220 ;
        RECT  4.540 0.505 6.890 0.735 ;
        RECT  5.985 0.965 6.215 2.785 ;
        RECT  4.585 0.965 5.985 1.195 ;
        RECT  5.725 2.555 5.985 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.415 0.965 4.585 1.250 ;
        RECT  3.575 1.020 4.415 1.250 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.590 0.465 2.960 ;
    END
END SEDFCND1BWP7T

MACRO SEDFCND2BWP7T
    CLASS CORE ;
    FOREIGN SEDFCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.840 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.160 0.465 19.505 2.535 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.885 1.055 21.140 2.690 ;
        RECT  20.860 0.465 20.885 3.310 ;
        RECT  20.650 0.465 20.860 1.285 ;
        RECT  20.655 2.460 20.860 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.820 8.340 2.115 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4014 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.985 3.190 15.715 3.420 ;
        RECT  14.755 2.730 14.985 3.420 ;
        RECT  13.790 2.730 14.755 2.960 ;
        RECT  13.560 2.730 13.790 3.270 ;
        RECT  11.785 2.940 13.560 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.605 -0.235 21.840 0.235 ;
        RECT  21.375 -0.235 21.605 1.245 ;
        RECT  20.220 -0.235 21.375 0.235 ;
        RECT  19.880 -0.235 20.220 1.180 ;
        RECT  18.740 -0.235 19.880 0.235 ;
        RECT  18.400 -0.235 18.740 0.465 ;
        RECT  16.810 -0.235 18.400 0.235 ;
        RECT  16.470 -0.235 16.810 0.465 ;
        RECT  12.815 -0.235 16.470 0.235 ;
        RECT  12.475 -0.235 12.815 0.730 ;
        RECT  8.670 -0.235 12.475 0.235 ;
        RECT  8.330 -0.235 8.670 0.465 ;
        RECT  4.035 -0.235 8.330 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.605 3.685 21.840 4.155 ;
        RECT  21.375 2.255 21.605 4.155 ;
        RECT  20.220 3.685 21.375 4.155 ;
        RECT  19.880 3.250 20.220 4.155 ;
        RECT  18.625 3.685 19.880 4.155 ;
        RECT  18.285 3.250 18.625 4.155 ;
        RECT  17.055 3.685 18.285 4.155 ;
        RECT  16.715 3.190 17.055 4.155 ;
        RECT  14.480 3.685 16.715 4.155 ;
        RECT  14.140 3.190 14.480 4.155 ;
        RECT  8.205 3.685 14.140 4.155 ;
        RECT  7.865 3.440 8.205 4.155 ;
        RECT  3.995 3.685 7.865 4.155 ;
        RECT  3.635 2.950 3.995 4.155 ;
        RECT  1.290 3.685 3.635 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  20.175 1.600 20.405 3.020 ;
        RECT  18.430 2.790 20.175 3.020 ;
        RECT  18.690 0.695 18.920 1.940 ;
        RECT  15.995 0.695 18.690 0.925 ;
        RECT  18.200 1.155 18.430 3.020 ;
        RECT  16.985 1.155 18.200 1.385 ;
        RECT  17.775 2.540 18.200 2.770 ;
        RECT  17.670 1.670 17.900 2.260 ;
        RECT  17.545 2.540 17.775 3.370 ;
        RECT  17.005 2.030 17.670 2.260 ;
        RECT  16.775 2.030 17.005 2.960 ;
        RECT  16.755 1.155 16.985 1.800 ;
        RECT  15.445 2.730 16.775 2.960 ;
        RECT  16.255 1.570 16.755 1.800 ;
        RECT  15.995 2.270 16.220 2.500 ;
        RECT  15.765 0.465 15.995 2.500 ;
        RECT  15.195 1.045 15.765 1.275 ;
        RECT  15.215 1.615 15.445 2.960 ;
        RECT  14.605 1.615 15.215 1.845 ;
        RECT  14.965 0.465 15.195 1.275 ;
        RECT  13.275 0.465 14.965 0.695 ;
        RECT  14.375 0.990 14.605 1.845 ;
        RECT  13.990 2.270 14.585 2.500 ;
        RECT  14.150 0.990 14.375 1.220 ;
        RECT  13.760 1.420 13.990 2.500 ;
        RECT  13.735 1.420 13.760 1.650 ;
        RECT  13.505 0.925 13.735 1.650 ;
        RECT  12.725 1.420 13.505 1.650 ;
        RECT  13.055 1.880 13.395 2.200 ;
        RECT  13.045 0.465 13.275 1.190 ;
        RECT  11.545 2.440 13.205 2.670 ;
        RECT  11.025 1.970 13.055 2.200 ;
        RECT  11.780 0.960 13.045 1.190 ;
        RECT  12.385 1.420 12.725 1.740 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  9.135 0.465 11.550 0.695 ;
        RECT  11.020 1.970 11.025 2.725 ;
        RECT  10.790 0.935 11.020 2.725 ;
        RECT  10.255 0.990 10.390 2.865 ;
        RECT  10.155 0.990 10.255 3.210 ;
        RECT  9.965 0.990 10.155 1.220 ;
        RECT  10.025 2.525 10.155 3.210 ;
        RECT  7.775 2.980 10.025 3.210 ;
        RECT  9.725 1.805 9.925 2.035 ;
        RECT  9.495 1.115 9.725 2.670 ;
        RECT  9.265 1.115 9.495 1.345 ;
        RECT  9.270 2.440 9.495 2.670 ;
        RECT  9.005 1.800 9.200 2.040 ;
        RECT  8.905 0.465 9.135 0.925 ;
        RECT  8.775 1.155 9.005 2.725 ;
        RECT  7.700 0.695 8.905 0.925 ;
        RECT  7.940 1.155 8.775 1.385 ;
        RECT  8.005 2.380 8.775 2.725 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.470 0.695 7.700 1.590 ;
        RECT  6.215 2.555 7.545 2.785 ;
        RECT  6.935 1.360 7.470 1.590 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.890 0.505 7.230 1.130 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  6.705 1.360 6.935 2.220 ;
        RECT  4.540 0.505 6.890 0.735 ;
        RECT  5.985 0.965 6.215 2.785 ;
        RECT  4.585 0.965 5.985 1.195 ;
        RECT  5.725 2.555 5.985 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.415 0.965 4.585 1.250 ;
        RECT  3.575 1.020 4.415 1.250 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.590 0.465 2.960 ;
    END
END SEDFCND2BWP7T

MACRO SEDFCNQD0BWP7T
    CLASS CORE ;
    FOREIGN SEDFCNQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.130 0.495 19.460 2.715 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.820 8.340 2.115 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4068 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.160 2.395 17.275 2.625 ;
        RECT  16.930 2.395 17.160 3.455 ;
        RECT  14.940 3.225 16.930 3.455 ;
        RECT  14.710 2.730 14.940 3.455 ;
        RECT  13.790 2.730 14.710 2.960 ;
        RECT  13.560 2.730 13.790 3.270 ;
        RECT  11.785 2.940 13.560 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.700 -0.235 19.600 0.235 ;
        RECT  18.360 -0.235 18.700 0.790 ;
        RECT  16.175 -0.235 18.360 0.235 ;
        RECT  15.835 -0.235 16.175 0.465 ;
        RECT  12.815 -0.235 15.835 0.235 ;
        RECT  12.475 -0.235 12.815 0.730 ;
        RECT  8.670 -0.235 12.475 0.235 ;
        RECT  8.330 -0.235 8.670 0.465 ;
        RECT  4.035 -0.235 8.330 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.615 3.685 19.600 4.155 ;
        RECT  18.275 2.850 18.615 4.155 ;
        RECT  14.480 3.685 18.275 4.155 ;
        RECT  14.140 3.190 14.480 4.155 ;
        RECT  8.205 3.685 14.140 4.155 ;
        RECT  7.865 3.440 8.205 4.155 ;
        RECT  3.995 3.685 7.865 4.155 ;
        RECT  3.635 2.950 3.995 4.155 ;
        RECT  1.290 3.685 3.635 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.580 1.600 18.885 1.940 ;
        RECT  18.350 1.020 18.580 2.620 ;
        RECT  17.945 1.020 18.350 1.250 ;
        RECT  17.740 2.390 18.350 2.620 ;
        RECT  17.725 1.565 17.955 2.160 ;
        RECT  17.715 0.495 17.945 1.250 ;
        RECT  17.510 2.390 17.740 3.200 ;
        RECT  16.700 1.930 17.725 2.160 ;
        RECT  17.070 1.020 17.715 1.250 ;
        RECT  16.840 1.020 17.070 1.700 ;
        RECT  16.090 1.470 16.840 1.700 ;
        RECT  16.470 1.930 16.700 2.995 ;
        RECT  15.400 2.765 16.470 2.995 ;
        RECT  15.860 0.950 16.190 1.180 ;
        RECT  15.860 2.305 16.190 2.535 ;
        RECT  15.630 0.950 15.860 2.535 ;
        RECT  15.165 0.950 15.630 1.220 ;
        RECT  15.170 1.615 15.400 2.995 ;
        RECT  14.610 1.615 15.170 1.845 ;
        RECT  14.935 0.465 15.165 1.220 ;
        RECT  13.275 0.465 14.935 0.695 ;
        RECT  14.380 0.990 14.610 1.845 ;
        RECT  13.990 2.270 14.505 2.500 ;
        RECT  14.150 0.990 14.380 1.220 ;
        RECT  13.760 1.420 13.990 2.500 ;
        RECT  13.735 1.420 13.760 1.650 ;
        RECT  13.505 0.925 13.735 1.650 ;
        RECT  12.725 1.420 13.505 1.650 ;
        RECT  13.055 1.880 13.395 2.200 ;
        RECT  13.045 0.465 13.275 1.190 ;
        RECT  11.545 2.440 13.205 2.670 ;
        RECT  11.025 1.970 13.055 2.200 ;
        RECT  11.780 0.960 13.045 1.190 ;
        RECT  12.385 1.420 12.725 1.740 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  9.135 0.465 11.550 0.695 ;
        RECT  11.020 1.970 11.025 2.725 ;
        RECT  10.790 0.935 11.020 2.725 ;
        RECT  10.255 0.990 10.390 2.865 ;
        RECT  10.155 0.990 10.255 3.210 ;
        RECT  9.965 0.990 10.155 1.220 ;
        RECT  10.025 2.525 10.155 3.210 ;
        RECT  7.775 2.980 10.025 3.210 ;
        RECT  9.725 1.805 9.925 2.035 ;
        RECT  9.495 1.115 9.725 2.670 ;
        RECT  9.265 1.115 9.495 1.345 ;
        RECT  9.270 2.440 9.495 2.670 ;
        RECT  9.005 1.800 9.200 2.040 ;
        RECT  8.905 0.465 9.135 0.925 ;
        RECT  8.775 1.155 9.005 2.725 ;
        RECT  7.700 0.695 8.905 0.925 ;
        RECT  7.940 1.155 8.775 1.385 ;
        RECT  8.005 2.380 8.775 2.725 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.470 0.695 7.700 1.590 ;
        RECT  6.215 2.555 7.545 2.785 ;
        RECT  6.935 1.360 7.470 1.590 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.890 0.505 7.230 1.130 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  6.705 1.360 6.935 2.220 ;
        RECT  4.540 0.505 6.890 0.735 ;
        RECT  5.985 0.965 6.215 2.785 ;
        RECT  4.585 0.965 5.985 1.195 ;
        RECT  5.725 2.555 5.985 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.415 0.965 4.585 1.250 ;
        RECT  3.575 1.020 4.415 1.250 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.590 0.465 2.960 ;
    END
END SEDFCNQD0BWP7T

MACRO SEDFCNQD1BWP7T
    CLASS CORE ;
    FOREIGN SEDFCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.130 0.470 19.460 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.820 8.340 2.115 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4068 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.160 2.395 17.275 2.625 ;
        RECT  16.930 2.395 17.160 3.455 ;
        RECT  14.940 3.225 16.930 3.455 ;
        RECT  14.710 2.730 14.940 3.455 ;
        RECT  13.790 2.730 14.710 2.960 ;
        RECT  13.560 2.730 13.790 3.270 ;
        RECT  11.785 2.940 13.560 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.700 -0.235 19.600 0.235 ;
        RECT  18.360 -0.235 18.700 0.790 ;
        RECT  16.090 -0.235 18.360 0.235 ;
        RECT  15.750 -0.235 16.090 0.465 ;
        RECT  12.815 -0.235 15.750 0.235 ;
        RECT  12.475 -0.235 12.815 0.730 ;
        RECT  8.670 -0.235 12.475 0.235 ;
        RECT  8.330 -0.235 8.670 0.465 ;
        RECT  4.035 -0.235 8.330 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.595 3.685 19.600 4.155 ;
        RECT  18.255 2.850 18.595 4.155 ;
        RECT  14.480 3.685 18.255 4.155 ;
        RECT  14.140 3.190 14.480 4.155 ;
        RECT  8.205 3.685 14.140 4.155 ;
        RECT  7.865 3.440 8.205 4.155 ;
        RECT  3.995 3.685 7.865 4.155 ;
        RECT  3.635 2.950 3.995 4.155 ;
        RECT  1.290 3.685 3.635 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.580 1.600 18.885 1.940 ;
        RECT  18.350 1.020 18.580 2.620 ;
        RECT  17.945 1.020 18.350 1.250 ;
        RECT  17.740 2.390 18.350 2.620 ;
        RECT  17.715 0.495 17.945 1.250 ;
        RECT  17.705 1.565 17.935 2.160 ;
        RECT  17.510 2.390 17.740 3.200 ;
        RECT  17.070 1.020 17.715 1.250 ;
        RECT  16.700 1.930 17.705 2.160 ;
        RECT  16.840 1.020 17.070 1.700 ;
        RECT  16.090 1.470 16.840 1.700 ;
        RECT  16.470 1.930 16.700 2.995 ;
        RECT  15.400 2.765 16.470 2.995 ;
        RECT  15.860 0.950 16.190 1.180 ;
        RECT  15.860 2.305 16.190 2.535 ;
        RECT  15.630 0.950 15.860 2.535 ;
        RECT  15.165 0.950 15.630 1.220 ;
        RECT  15.170 1.615 15.400 2.995 ;
        RECT  14.610 1.615 15.170 1.845 ;
        RECT  14.935 0.465 15.165 1.220 ;
        RECT  13.275 0.465 14.935 0.695 ;
        RECT  14.380 0.990 14.610 1.845 ;
        RECT  13.990 2.270 14.505 2.500 ;
        RECT  14.150 0.990 14.380 1.220 ;
        RECT  13.760 1.420 13.990 2.500 ;
        RECT  13.735 1.420 13.760 1.650 ;
        RECT  13.505 0.925 13.735 1.650 ;
        RECT  12.725 1.420 13.505 1.650 ;
        RECT  13.055 1.880 13.395 2.200 ;
        RECT  13.045 0.465 13.275 1.190 ;
        RECT  11.545 2.440 13.205 2.670 ;
        RECT  11.025 1.970 13.055 2.200 ;
        RECT  11.780 0.960 13.045 1.190 ;
        RECT  12.385 1.420 12.725 1.740 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  9.135 0.465 11.550 0.695 ;
        RECT  11.020 1.970 11.025 2.725 ;
        RECT  10.790 0.935 11.020 2.725 ;
        RECT  10.255 0.990 10.390 2.865 ;
        RECT  10.155 0.990 10.255 3.210 ;
        RECT  9.965 0.990 10.155 1.220 ;
        RECT  10.025 2.525 10.155 3.210 ;
        RECT  7.775 2.980 10.025 3.210 ;
        RECT  9.725 1.805 9.925 2.035 ;
        RECT  9.495 1.115 9.725 2.670 ;
        RECT  9.265 1.115 9.495 1.345 ;
        RECT  9.270 2.440 9.495 2.670 ;
        RECT  9.005 1.800 9.200 2.040 ;
        RECT  8.905 0.465 9.135 0.925 ;
        RECT  8.775 1.155 9.005 2.725 ;
        RECT  7.700 0.695 8.905 0.925 ;
        RECT  7.940 1.155 8.775 1.385 ;
        RECT  8.005 2.380 8.775 2.725 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.470 0.695 7.700 1.590 ;
        RECT  6.215 2.555 7.545 2.785 ;
        RECT  6.935 1.360 7.470 1.590 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.890 0.505 7.230 1.130 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  6.705 1.360 6.935 2.220 ;
        RECT  4.540 0.505 6.890 0.735 ;
        RECT  5.985 0.965 6.215 2.785 ;
        RECT  4.585 0.965 5.985 1.195 ;
        RECT  5.725 2.555 5.985 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.415 0.965 4.585 1.250 ;
        RECT  3.575 1.020 4.415 1.250 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.590 0.465 2.960 ;
    END
END SEDFCNQD1BWP7T

MACRO SEDFCNQD2BWP7T
    CLASS CORE ;
    FOREIGN SEDFCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.205 1.060 19.460 2.730 ;
        RECT  19.180 0.470 19.205 3.310 ;
        RECT  18.975 0.470 19.180 1.290 ;
        RECT  18.975 2.495 19.180 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 1.820 8.340 2.115 ;
        END
    END CP
    PIN CDN
        ANTENNAGATEAREA 0.4068 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.160 2.395 17.275 2.625 ;
        RECT  16.930 2.395 17.160 3.455 ;
        RECT  14.940 3.225 16.930 3.455 ;
        RECT  14.710 2.730 14.940 3.455 ;
        RECT  13.790 2.730 14.710 2.960 ;
        RECT  13.560 2.730 13.790 3.270 ;
        RECT  11.785 2.940 13.560 3.270 ;
        END
    END CDN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.925 -0.235 20.160 0.235 ;
        RECT  19.695 -0.235 19.925 1.255 ;
        RECT  18.500 -0.235 19.695 0.235 ;
        RECT  18.160 -0.235 18.500 0.465 ;
        RECT  16.090 -0.235 18.160 0.235 ;
        RECT  15.750 -0.235 16.090 0.465 ;
        RECT  12.815 -0.235 15.750 0.235 ;
        RECT  12.475 -0.235 12.815 0.730 ;
        RECT  8.670 -0.235 12.475 0.235 ;
        RECT  8.330 -0.235 8.670 0.465 ;
        RECT  4.035 -0.235 8.330 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.925 3.685 20.160 4.155 ;
        RECT  19.695 2.250 19.925 4.155 ;
        RECT  18.535 3.685 19.695 4.155 ;
        RECT  18.195 2.940 18.535 4.155 ;
        RECT  14.480 3.685 18.195 4.155 ;
        RECT  14.140 3.190 14.480 4.155 ;
        RECT  8.205 3.685 14.140 4.155 ;
        RECT  7.865 3.440 8.205 4.155 ;
        RECT  3.995 3.685 7.865 4.155 ;
        RECT  3.635 2.950 3.995 4.155 ;
        RECT  1.290 3.685 3.635 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.435 1.020 18.665 2.620 ;
        RECT  17.070 1.020 18.435 1.250 ;
        RECT  17.740 2.390 18.435 2.620 ;
        RECT  17.675 1.565 17.905 2.160 ;
        RECT  17.510 2.390 17.740 3.200 ;
        RECT  16.675 1.930 17.675 2.160 ;
        RECT  16.840 1.020 17.070 1.700 ;
        RECT  16.090 1.470 16.840 1.700 ;
        RECT  16.445 1.930 16.675 2.995 ;
        RECT  15.400 2.765 16.445 2.995 ;
        RECT  15.860 2.305 16.190 2.535 ;
        RECT  15.860 0.950 16.140 1.180 ;
        RECT  15.630 0.950 15.860 2.535 ;
        RECT  15.165 0.950 15.630 1.220 ;
        RECT  15.170 1.615 15.400 2.995 ;
        RECT  14.610 1.615 15.170 1.845 ;
        RECT  14.935 0.465 15.165 1.220 ;
        RECT  13.275 0.465 14.935 0.695 ;
        RECT  14.380 0.990 14.610 1.845 ;
        RECT  13.990 2.270 14.505 2.500 ;
        RECT  14.150 0.990 14.380 1.220 ;
        RECT  13.760 1.420 13.990 2.500 ;
        RECT  13.735 1.420 13.760 1.650 ;
        RECT  13.505 0.925 13.735 1.650 ;
        RECT  12.725 1.420 13.505 1.650 ;
        RECT  13.055 1.880 13.395 2.200 ;
        RECT  13.045 0.465 13.275 1.190 ;
        RECT  11.545 2.440 13.205 2.670 ;
        RECT  11.025 1.970 13.055 2.200 ;
        RECT  11.780 0.960 13.045 1.190 ;
        RECT  12.385 1.420 12.725 1.740 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  9.135 0.465 11.550 0.695 ;
        RECT  11.020 1.970 11.025 2.725 ;
        RECT  10.790 0.935 11.020 2.725 ;
        RECT  10.255 0.990 10.390 2.865 ;
        RECT  10.155 0.990 10.255 3.210 ;
        RECT  9.965 0.990 10.155 1.220 ;
        RECT  10.025 2.525 10.155 3.210 ;
        RECT  7.775 2.980 10.025 3.210 ;
        RECT  9.725 1.805 9.925 2.035 ;
        RECT  9.495 1.115 9.725 2.670 ;
        RECT  9.265 1.115 9.495 1.345 ;
        RECT  9.270 2.440 9.495 2.670 ;
        RECT  9.005 1.800 9.200 2.040 ;
        RECT  8.905 0.465 9.135 0.925 ;
        RECT  8.775 1.155 9.005 2.725 ;
        RECT  7.700 0.695 8.905 0.925 ;
        RECT  7.940 1.155 8.775 1.385 ;
        RECT  8.005 2.380 8.775 2.725 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.470 0.695 7.700 1.590 ;
        RECT  6.215 2.555 7.545 2.785 ;
        RECT  6.935 1.360 7.470 1.590 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.890 0.505 7.230 1.130 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  6.705 1.360 6.935 2.220 ;
        RECT  4.540 0.505 6.890 0.735 ;
        RECT  5.985 0.965 6.215 2.785 ;
        RECT  4.585 0.965 5.985 1.195 ;
        RECT  5.725 2.555 5.985 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.415 0.965 4.585 1.250 ;
        RECT  3.575 1.020 4.415 1.250 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.590 0.465 2.960 ;
    END
END SEDFCNQD2BWP7T

MACRO SEDFD0BWP7T
    CLASS CORE ;
    FOREIGN SEDFD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.500 1.075 17.780 2.560 ;
        RECT  17.365 1.075 17.500 1.305 ;
        RECT  17.080 2.330 17.500 2.560 ;
        RECT  17.135 0.480 17.365 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.570 0.470 18.900 2.715 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.140 -0.235 19.040 0.235 ;
        RECT  17.800 -0.235 18.140 0.775 ;
        RECT  15.010 -0.235 17.800 0.235 ;
        RECT  14.780 -0.235 15.010 0.520 ;
        RECT  12.445 -0.235 14.780 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.075 3.685 19.040 4.155 ;
        RECT  17.735 3.340 18.075 4.155 ;
        RECT  15.940 3.685 17.735 4.155 ;
        RECT  15.595 3.225 15.940 4.155 ;
        RECT  12.600 3.685 15.595 4.155 ;
        RECT  12.240 3.190 12.600 4.155 ;
        RECT  8.905 3.685 12.240 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.095 1.600 18.325 3.020 ;
        RECT  16.850 2.790 18.095 3.020 ;
        RECT  15.470 0.465 16.900 0.695 ;
        RECT  16.660 1.020 16.850 3.020 ;
        RECT  16.620 1.020 16.660 3.380 ;
        RECT  15.930 1.020 16.620 1.250 ;
        RECT  16.430 2.790 16.620 3.380 ;
        RECT  16.160 1.595 16.390 2.455 ;
        RECT  15.855 2.225 16.160 2.455 ;
        RECT  15.700 1.020 15.930 1.885 ;
        RECT  15.625 2.225 15.855 2.995 ;
        RECT  15.010 1.655 15.700 1.885 ;
        RECT  14.090 2.765 15.625 2.995 ;
        RECT  15.240 0.465 15.470 1.220 ;
        RECT  14.550 0.990 15.240 1.220 ;
        RECT  14.550 2.300 15.085 2.530 ;
        RECT  13.350 3.225 14.750 3.455 ;
        RECT  14.320 0.465 14.550 2.530 ;
        RECT  12.905 0.465 14.320 0.695 ;
        RECT  13.860 0.925 14.090 2.995 ;
        RECT  13.365 1.420 13.505 2.500 ;
        RECT  13.275 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  13.135 0.925 13.275 1.650 ;
        RECT  13.085 2.270 13.275 2.500 ;
        RECT  12.175 1.420 13.135 1.650 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.515 1.880 12.855 2.415 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  11.200 2.185 12.515 2.415 ;
        RECT  11.835 1.420 12.175 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFD0BWP7T

MACRO SEDFD1BWP7T
    CLASS CORE ;
    FOREIGN SEDFD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.500 1.075 17.780 2.560 ;
        RECT  17.365 1.075 17.500 1.305 ;
        RECT  17.080 2.330 17.500 2.560 ;
        RECT  17.135 0.480 17.365 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.570 0.470 18.900 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.140 -0.235 19.040 0.235 ;
        RECT  17.800 -0.235 18.140 0.810 ;
        RECT  15.010 -0.235 17.800 0.235 ;
        RECT  14.780 -0.235 15.010 0.520 ;
        RECT  12.445 -0.235 14.780 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.140 3.685 19.040 4.155 ;
        RECT  17.800 3.250 18.140 4.155 ;
        RECT  15.995 3.685 17.800 4.155 ;
        RECT  15.650 3.225 15.995 4.155 ;
        RECT  12.600 3.685 15.650 4.155 ;
        RECT  12.240 3.190 12.600 4.155 ;
        RECT  8.905 3.685 12.240 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.095 1.600 18.325 3.020 ;
        RECT  16.850 2.790 18.095 3.020 ;
        RECT  15.470 0.465 16.900 0.695 ;
        RECT  16.660 1.020 16.850 3.020 ;
        RECT  16.620 1.020 16.660 3.380 ;
        RECT  15.930 1.020 16.620 1.250 ;
        RECT  16.430 2.565 16.620 3.380 ;
        RECT  16.160 1.530 16.390 2.300 ;
        RECT  15.855 2.070 16.160 2.300 ;
        RECT  15.700 1.020 15.930 1.830 ;
        RECT  15.625 2.070 15.855 2.995 ;
        RECT  15.010 1.600 15.700 1.830 ;
        RECT  14.090 2.765 15.625 2.995 ;
        RECT  15.240 0.465 15.470 1.220 ;
        RECT  14.550 0.990 15.240 1.220 ;
        RECT  14.550 2.300 15.085 2.530 ;
        RECT  13.350 3.225 14.750 3.455 ;
        RECT  14.320 0.465 14.550 2.530 ;
        RECT  12.905 0.465 14.320 0.695 ;
        RECT  13.860 0.925 14.090 2.995 ;
        RECT  13.365 1.420 13.505 2.500 ;
        RECT  13.275 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  13.135 0.925 13.275 1.650 ;
        RECT  13.085 2.270 13.275 2.500 ;
        RECT  12.175 1.420 13.135 1.650 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.515 1.880 12.855 2.415 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  11.200 2.185 12.515 2.415 ;
        RECT  11.835 1.420 12.175 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFD1BWP7T

MACRO SEDFD2BWP7T
    CLASS CORE ;
    FOREIGN SEDFD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3206 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.480 0.495 17.820 2.530 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.205 1.060 19.460 2.735 ;
        RECT  19.180 0.480 19.205 3.310 ;
        RECT  18.975 0.480 19.180 1.290 ;
        RECT  18.975 2.500 19.180 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.925 -0.235 20.160 0.235 ;
        RECT  19.695 -0.235 19.925 1.275 ;
        RECT  18.540 -0.235 19.695 0.235 ;
        RECT  18.200 -0.235 18.540 0.810 ;
        RECT  17.060 -0.235 18.200 0.235 ;
        RECT  16.720 -0.235 17.060 0.465 ;
        RECT  15.760 -0.235 16.720 0.235 ;
        RECT  15.420 -0.235 15.760 0.465 ;
        RECT  12.445 -0.235 15.420 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.925 3.685 20.160 4.155 ;
        RECT  19.695 2.255 19.925 4.155 ;
        RECT  18.540 3.685 19.695 4.155 ;
        RECT  18.200 3.250 18.540 4.155 ;
        RECT  17.060 3.685 18.200 4.155 ;
        RECT  16.720 3.250 17.060 4.155 ;
        RECT  15.630 3.685 16.720 4.155 ;
        RECT  15.285 3.225 15.630 4.155 ;
        RECT  12.600 3.685 15.285 4.155 ;
        RECT  12.240 3.190 12.600 4.155 ;
        RECT  8.905 3.685 12.240 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.495 1.600 18.725 3.020 ;
        RECT  16.625 2.790 18.495 3.020 ;
        RECT  16.925 0.695 17.155 1.940 ;
        RECT  14.895 0.695 16.925 0.925 ;
        RECT  16.395 1.155 16.625 3.020 ;
        RECT  15.545 1.155 16.395 1.385 ;
        RECT  16.295 2.565 16.395 3.020 ;
        RECT  16.065 2.565 16.295 3.380 ;
        RECT  15.880 1.695 16.110 2.300 ;
        RECT  15.540 2.070 15.880 2.300 ;
        RECT  15.315 1.155 15.545 1.840 ;
        RECT  15.310 2.070 15.540 2.995 ;
        RECT  14.870 1.610 15.315 1.840 ;
        RECT  14.090 2.765 15.310 2.995 ;
        RECT  14.665 0.465 14.895 1.380 ;
        RECT  14.580 2.300 14.870 2.530 ;
        RECT  12.905 0.465 14.665 0.695 ;
        RECT  14.580 1.150 14.665 1.380 ;
        RECT  14.350 1.150 14.580 2.530 ;
        RECT  13.350 3.225 14.480 3.455 ;
        RECT  13.825 0.935 14.090 2.995 ;
        RECT  13.365 1.420 13.505 2.500 ;
        RECT  13.275 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  13.135 0.925 13.275 1.650 ;
        RECT  13.050 2.270 13.275 2.500 ;
        RECT  12.165 1.420 13.135 1.650 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.640 1.880 12.835 2.110 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  12.410 1.880 12.640 2.415 ;
        RECT  11.200 2.185 12.410 2.415 ;
        RECT  11.825 1.420 12.165 1.875 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFD2BWP7T

MACRO SEDFKCND0BWP7T
    CLASS CORE ;
    FOREIGN SEDFKCND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.620 1.075 18.900 2.560 ;
        RECT  18.485 1.075 18.620 1.305 ;
        RECT  18.200 2.330 18.620 2.560 ;
        RECT  18.255 0.480 18.485 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.690 0.470 20.020 2.715 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4581 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.820 6.630 2.100 ;
        RECT  5.380 1.540 5.720 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.765 9.940 2.710 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1782 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 2.370 6.860 2.660 ;
        RECT  4.755 1.485 4.985 2.660 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.260 -0.235 20.160 0.235 ;
        RECT  18.920 -0.235 19.260 0.775 ;
        RECT  16.130 -0.235 18.920 0.235 ;
        RECT  15.900 -0.235 16.130 0.520 ;
        RECT  13.565 -0.235 15.900 0.235 ;
        RECT  13.225 -0.235 13.565 0.730 ;
        RECT  9.845 -0.235 13.225 0.235 ;
        RECT  9.505 -0.235 9.845 0.465 ;
        RECT  4.035 -0.235 9.505 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.195 3.685 20.160 4.155 ;
        RECT  18.855 3.340 19.195 4.155 ;
        RECT  17.060 3.685 18.855 4.155 ;
        RECT  16.715 3.225 17.060 4.155 ;
        RECT  13.720 3.685 16.715 4.155 ;
        RECT  13.360 3.190 13.720 4.155 ;
        RECT  10.025 3.685 13.360 4.155 ;
        RECT  9.685 3.455 10.025 4.155 ;
        RECT  3.940 3.685 9.685 4.155 ;
        RECT  3.580 2.960 3.940 4.155 ;
        RECT  1.290 3.685 3.580 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.215 1.600 19.445 3.020 ;
        RECT  17.970 2.790 19.215 3.020 ;
        RECT  16.590 0.465 18.020 0.695 ;
        RECT  17.780 1.020 17.970 3.020 ;
        RECT  17.740 1.020 17.780 3.380 ;
        RECT  17.050 1.020 17.740 1.250 ;
        RECT  17.550 2.790 17.740 3.380 ;
        RECT  17.280 1.595 17.510 2.455 ;
        RECT  16.975 2.225 17.280 2.455 ;
        RECT  16.820 1.020 17.050 1.885 ;
        RECT  16.745 2.225 16.975 2.995 ;
        RECT  16.130 1.655 16.820 1.885 ;
        RECT  15.210 2.765 16.745 2.995 ;
        RECT  16.360 0.465 16.590 1.220 ;
        RECT  15.670 0.990 16.360 1.220 ;
        RECT  15.670 2.300 16.205 2.530 ;
        RECT  14.470 3.225 15.870 3.455 ;
        RECT  15.440 0.465 15.670 2.530 ;
        RECT  14.025 0.465 15.440 0.695 ;
        RECT  14.980 0.925 15.210 2.995 ;
        RECT  14.485 1.420 14.625 2.500 ;
        RECT  14.395 0.925 14.485 2.500 ;
        RECT  14.240 2.730 14.470 3.455 ;
        RECT  14.255 0.925 14.395 1.650 ;
        RECT  14.205 2.270 14.395 2.500 ;
        RECT  13.295 1.420 14.255 1.650 ;
        RECT  12.955 2.730 14.240 2.960 ;
        RECT  13.795 0.465 14.025 1.190 ;
        RECT  13.635 1.880 13.975 2.415 ;
        RECT  12.900 0.960 13.795 1.190 ;
        RECT  12.320 2.185 13.635 2.415 ;
        RECT  12.955 1.420 13.295 1.835 ;
        RECT  12.725 2.730 12.955 3.250 ;
        RECT  12.670 0.465 12.900 1.190 ;
        RECT  11.755 3.020 12.725 3.250 ;
        RECT  10.350 0.465 12.670 0.695 ;
        RECT  12.090 0.935 12.320 2.705 ;
        RECT  11.525 0.925 11.755 2.585 ;
        RECT  11.310 0.925 11.525 1.155 ;
        RECT  11.295 2.345 11.525 3.210 ;
        RECT  11.035 1.615 11.295 1.955 ;
        RECT  8.945 2.980 11.295 3.210 ;
        RECT  10.805 0.925 11.035 2.750 ;
        RECT  10.670 0.925 10.805 1.265 ;
        RECT  10.515 2.520 10.805 2.750 ;
        RECT  10.420 1.770 10.560 2.110 ;
        RECT  10.190 1.155 10.420 2.110 ;
        RECT  10.120 0.465 10.350 0.925 ;
        RECT  9.405 1.155 10.190 1.385 ;
        RECT  8.555 0.695 10.120 0.925 ;
        RECT  9.175 1.155 9.405 2.750 ;
        RECT  8.865 1.155 9.175 1.385 ;
        RECT  8.715 2.120 8.945 3.210 ;
        RECT  7.335 2.120 8.715 2.350 ;
        RECT  8.325 0.695 8.555 1.860 ;
        RECT  8.255 2.645 8.485 3.455 ;
        RECT  7.565 1.630 8.325 1.860 ;
        RECT  6.630 3.225 8.255 3.455 ;
        RECT  7.825 0.505 8.055 1.315 ;
        RECT  5.095 0.505 7.825 0.735 ;
        RECT  7.105 1.020 7.335 2.985 ;
        RECT  3.575 1.020 7.105 1.250 ;
        RECT  6.290 2.910 6.630 3.455 ;
        RECT  4.730 3.225 6.290 3.455 ;
        RECT  4.390 2.960 4.730 3.455 ;
        RECT  4.020 1.480 4.375 1.770 ;
        RECT  3.115 1.480 4.020 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFKCND0BWP7T

MACRO SEDFKCND1BWP7T
    CLASS CORE ;
    FOREIGN SEDFKCND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.160 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1088 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.620 1.075 18.900 2.560 ;
        RECT  18.485 1.075 18.620 1.305 ;
        RECT  18.200 2.330 18.620 2.560 ;
        RECT  18.255 0.480 18.485 1.305 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.690 0.470 20.020 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4581 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.820 6.630 2.100 ;
        RECT  5.380 1.540 5.720 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.765 9.940 2.710 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1782 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 2.370 6.860 2.660 ;
        RECT  4.755 1.485 4.985 2.660 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.260 -0.235 20.160 0.235 ;
        RECT  18.920 -0.235 19.260 0.810 ;
        RECT  16.130 -0.235 18.920 0.235 ;
        RECT  15.900 -0.235 16.130 0.520 ;
        RECT  13.565 -0.235 15.900 0.235 ;
        RECT  13.225 -0.235 13.565 0.730 ;
        RECT  9.845 -0.235 13.225 0.235 ;
        RECT  9.505 -0.235 9.845 0.465 ;
        RECT  4.035 -0.235 9.505 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.260 3.685 20.160 4.155 ;
        RECT  18.920 3.250 19.260 4.155 ;
        RECT  17.115 3.685 18.920 4.155 ;
        RECT  16.770 3.225 17.115 4.155 ;
        RECT  13.720 3.685 16.770 4.155 ;
        RECT  13.360 3.190 13.720 4.155 ;
        RECT  10.025 3.685 13.360 4.155 ;
        RECT  9.685 3.455 10.025 4.155 ;
        RECT  3.940 3.685 9.685 4.155 ;
        RECT  3.580 2.960 3.940 4.155 ;
        RECT  1.290 3.685 3.580 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.215 1.600 19.445 3.020 ;
        RECT  17.970 2.790 19.215 3.020 ;
        RECT  16.590 0.465 18.020 0.695 ;
        RECT  17.780 1.020 17.970 3.020 ;
        RECT  17.740 1.020 17.780 3.380 ;
        RECT  17.050 1.020 17.740 1.250 ;
        RECT  17.550 2.565 17.740 3.380 ;
        RECT  17.280 1.530 17.510 2.300 ;
        RECT  16.975 2.070 17.280 2.300 ;
        RECT  16.820 1.020 17.050 1.830 ;
        RECT  16.745 2.070 16.975 2.995 ;
        RECT  16.130 1.600 16.820 1.830 ;
        RECT  15.210 2.765 16.745 2.995 ;
        RECT  16.360 0.465 16.590 1.220 ;
        RECT  15.670 0.990 16.360 1.220 ;
        RECT  15.670 2.300 16.205 2.530 ;
        RECT  14.470 3.225 15.870 3.455 ;
        RECT  15.440 0.465 15.670 2.530 ;
        RECT  14.025 0.465 15.440 0.695 ;
        RECT  14.980 0.925 15.210 2.995 ;
        RECT  14.485 1.420 14.625 2.500 ;
        RECT  14.395 0.925 14.485 2.500 ;
        RECT  14.240 2.730 14.470 3.455 ;
        RECT  14.255 0.925 14.395 1.650 ;
        RECT  14.205 2.270 14.395 2.500 ;
        RECT  13.295 1.420 14.255 1.650 ;
        RECT  12.955 2.730 14.240 2.960 ;
        RECT  13.795 0.465 14.025 1.190 ;
        RECT  13.635 1.880 13.975 2.415 ;
        RECT  12.900 0.960 13.795 1.190 ;
        RECT  12.320 2.185 13.635 2.415 ;
        RECT  12.955 1.420 13.295 1.835 ;
        RECT  12.725 2.730 12.955 3.250 ;
        RECT  12.670 0.465 12.900 1.190 ;
        RECT  11.755 3.020 12.725 3.250 ;
        RECT  10.350 0.465 12.670 0.695 ;
        RECT  12.090 0.935 12.320 2.705 ;
        RECT  11.525 0.925 11.755 2.585 ;
        RECT  11.310 0.925 11.525 1.155 ;
        RECT  11.295 2.345 11.525 3.210 ;
        RECT  11.035 1.615 11.295 1.955 ;
        RECT  8.945 2.980 11.295 3.210 ;
        RECT  10.805 0.925 11.035 2.750 ;
        RECT  10.670 0.925 10.805 1.265 ;
        RECT  10.515 2.520 10.805 2.750 ;
        RECT  10.420 1.770 10.560 2.110 ;
        RECT  10.190 1.155 10.420 2.110 ;
        RECT  10.120 0.465 10.350 0.925 ;
        RECT  9.405 1.155 10.190 1.385 ;
        RECT  8.555 0.695 10.120 0.925 ;
        RECT  9.175 1.155 9.405 2.750 ;
        RECT  8.865 1.155 9.175 1.385 ;
        RECT  8.715 2.120 8.945 3.210 ;
        RECT  7.335 2.120 8.715 2.350 ;
        RECT  8.325 0.695 8.555 1.860 ;
        RECT  8.255 2.645 8.485 3.455 ;
        RECT  7.565 1.630 8.325 1.860 ;
        RECT  6.630 3.225 8.255 3.455 ;
        RECT  7.825 0.505 8.055 1.315 ;
        RECT  5.095 0.505 7.825 0.735 ;
        RECT  7.105 1.020 7.335 2.985 ;
        RECT  3.575 1.020 7.105 1.250 ;
        RECT  6.290 2.910 6.630 3.455 ;
        RECT  4.730 3.225 6.290 3.455 ;
        RECT  4.390 2.960 4.730 3.455 ;
        RECT  4.020 1.480 4.375 1.770 ;
        RECT  3.115 1.480 4.020 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFKCND1BWP7T

MACRO SEDFKCND2BWP7T
    CLASS CORE ;
    FOREIGN SEDFKCND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 21.280 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.3211 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.600 0.495 18.940 2.530 ;
        END
    END QN
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.325 1.060 20.580 2.735 ;
        RECT  20.300 0.480 20.325 3.310 ;
        RECT  20.095 0.480 20.300 1.290 ;
        RECT  20.095 2.500 20.300 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4581 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.820 6.630 2.100 ;
        RECT  5.380 1.540 5.720 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.765 9.940 2.710 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1782 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 2.370 6.860 2.660 ;
        RECT  4.755 1.485 4.985 2.660 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.045 -0.235 21.280 0.235 ;
        RECT  20.815 -0.235 21.045 1.275 ;
        RECT  19.660 -0.235 20.815 0.235 ;
        RECT  19.320 -0.235 19.660 0.810 ;
        RECT  18.180 -0.235 19.320 0.235 ;
        RECT  17.840 -0.235 18.180 0.465 ;
        RECT  16.880 -0.235 17.840 0.235 ;
        RECT  16.540 -0.235 16.880 0.465 ;
        RECT  13.565 -0.235 16.540 0.235 ;
        RECT  13.225 -0.235 13.565 0.730 ;
        RECT  9.845 -0.235 13.225 0.235 ;
        RECT  9.505 -0.235 9.845 0.465 ;
        RECT  4.035 -0.235 9.505 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.045 3.685 21.280 4.155 ;
        RECT  20.815 2.255 21.045 4.155 ;
        RECT  19.660 3.685 20.815 4.155 ;
        RECT  19.320 3.250 19.660 4.155 ;
        RECT  18.180 3.685 19.320 4.155 ;
        RECT  17.840 3.250 18.180 4.155 ;
        RECT  16.750 3.685 17.840 4.155 ;
        RECT  16.405 3.225 16.750 4.155 ;
        RECT  13.720 3.685 16.405 4.155 ;
        RECT  13.360 3.190 13.720 4.155 ;
        RECT  10.025 3.685 13.360 4.155 ;
        RECT  9.685 3.455 10.025 4.155 ;
        RECT  3.940 3.685 9.685 4.155 ;
        RECT  3.580 2.960 3.940 4.155 ;
        RECT  1.290 3.685 3.580 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.615 1.600 19.845 3.020 ;
        RECT  17.745 2.790 19.615 3.020 ;
        RECT  18.045 0.695 18.275 1.940 ;
        RECT  16.015 0.695 18.045 0.925 ;
        RECT  17.515 1.155 17.745 3.020 ;
        RECT  16.665 1.155 17.515 1.385 ;
        RECT  17.415 2.565 17.515 3.020 ;
        RECT  17.185 2.565 17.415 3.380 ;
        RECT  17.000 1.695 17.230 2.300 ;
        RECT  16.660 2.070 17.000 2.300 ;
        RECT  16.435 1.155 16.665 1.840 ;
        RECT  16.430 2.070 16.660 2.995 ;
        RECT  15.990 1.610 16.435 1.840 ;
        RECT  15.210 2.765 16.430 2.995 ;
        RECT  15.785 0.465 16.015 1.380 ;
        RECT  15.700 2.300 16.005 2.530 ;
        RECT  14.025 0.465 15.785 0.695 ;
        RECT  15.700 1.150 15.785 1.380 ;
        RECT  15.470 1.150 15.700 2.530 ;
        RECT  14.470 3.225 15.615 3.455 ;
        RECT  14.960 0.935 15.210 2.995 ;
        RECT  14.485 1.420 14.625 2.500 ;
        RECT  14.395 0.925 14.485 2.500 ;
        RECT  14.240 2.730 14.470 3.455 ;
        RECT  14.255 0.925 14.395 1.650 ;
        RECT  14.185 2.270 14.395 2.500 ;
        RECT  13.285 1.420 14.255 1.650 ;
        RECT  12.955 2.730 14.240 2.960 ;
        RECT  13.795 0.465 14.025 1.190 ;
        RECT  13.615 1.880 13.955 2.415 ;
        RECT  12.900 0.960 13.795 1.190 ;
        RECT  12.320 2.185 13.615 2.415 ;
        RECT  12.945 1.420 13.285 1.835 ;
        RECT  12.725 2.730 12.955 3.250 ;
        RECT  12.670 0.465 12.900 1.190 ;
        RECT  11.755 3.020 12.725 3.250 ;
        RECT  10.350 0.465 12.670 0.695 ;
        RECT  12.090 0.935 12.320 2.705 ;
        RECT  11.525 0.925 11.755 2.585 ;
        RECT  11.310 0.925 11.525 1.155 ;
        RECT  11.295 2.345 11.525 3.210 ;
        RECT  11.035 1.615 11.295 1.955 ;
        RECT  8.945 2.980 11.295 3.210 ;
        RECT  10.805 0.925 11.035 2.750 ;
        RECT  10.670 0.925 10.805 1.265 ;
        RECT  10.515 2.520 10.805 2.750 ;
        RECT  10.420 1.770 10.560 2.110 ;
        RECT  10.190 1.155 10.420 2.110 ;
        RECT  10.120 0.465 10.350 0.925 ;
        RECT  9.405 1.155 10.190 1.385 ;
        RECT  8.555 0.695 10.120 0.925 ;
        RECT  9.175 1.155 9.405 2.750 ;
        RECT  8.865 1.155 9.175 1.385 ;
        RECT  8.715 2.120 8.945 3.210 ;
        RECT  7.335 2.120 8.715 2.350 ;
        RECT  8.325 0.695 8.555 1.860 ;
        RECT  8.255 2.645 8.485 3.455 ;
        RECT  7.565 1.630 8.325 1.860 ;
        RECT  6.630 3.225 8.255 3.455 ;
        RECT  7.825 0.505 8.055 1.315 ;
        RECT  5.095 0.505 7.825 0.735 ;
        RECT  7.105 1.020 7.335 2.985 ;
        RECT  3.575 1.020 7.105 1.250 ;
        RECT  6.290 2.910 6.630 3.455 ;
        RECT  4.730 3.225 6.290 3.455 ;
        RECT  4.390 2.960 4.730 3.455 ;
        RECT  4.020 1.480 4.375 1.770 ;
        RECT  3.115 1.480 4.020 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFKCND2BWP7T

MACRO SEDFKCNQD0BWP7T
    CLASS CORE ;
    FOREIGN SEDFKCNQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.570 0.505 18.900 3.185 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4581 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.820 6.630 2.100 ;
        RECT  5.380 1.540 5.720 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.765 9.940 2.710 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1782 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 2.370 6.860 2.660 ;
        RECT  4.755 1.485 4.985 2.660 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.085 -0.235 19.040 0.235 ;
        RECT  17.855 -0.235 18.085 0.855 ;
        RECT  16.665 -0.235 17.855 0.235 ;
        RECT  16.325 -0.235 16.665 0.465 ;
        RECT  13.565 -0.235 16.325 0.235 ;
        RECT  13.225 -0.235 13.565 0.730 ;
        RECT  9.845 -0.235 13.225 0.235 ;
        RECT  9.505 -0.235 9.845 0.465 ;
        RECT  4.035 -0.235 9.505 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.085 3.685 19.040 4.155 ;
        RECT  17.855 2.850 18.085 4.155 ;
        RECT  16.680 3.685 17.855 4.155 ;
        RECT  16.340 3.455 16.680 4.155 ;
        RECT  13.720 3.685 16.340 4.155 ;
        RECT  13.360 3.190 13.720 4.155 ;
        RECT  10.025 3.685 13.360 4.155 ;
        RECT  9.685 3.455 10.025 4.155 ;
        RECT  3.940 3.685 9.685 4.155 ;
        RECT  3.580 2.960 3.940 4.155 ;
        RECT  1.290 3.685 3.580 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.620 1.600 18.325 1.940 ;
        RECT  17.390 0.960 17.620 2.750 ;
        RECT  16.635 0.960 17.390 1.190 ;
        RECT  17.100 2.520 17.390 2.750 ;
        RECT  16.930 1.565 17.160 2.290 ;
        RECT  16.730 2.060 16.930 2.290 ;
        RECT  16.500 2.060 16.730 2.995 ;
        RECT  16.405 0.960 16.635 1.830 ;
        RECT  15.210 2.765 16.500 2.995 ;
        RECT  16.120 1.600 16.405 1.830 ;
        RECT  15.810 2.300 16.135 2.530 ;
        RECT  15.810 0.990 16.120 1.220 ;
        RECT  14.470 3.225 15.845 3.455 ;
        RECT  15.580 0.465 15.810 2.530 ;
        RECT  14.025 0.465 15.580 0.695 ;
        RECT  14.980 0.925 15.210 2.995 ;
        RECT  14.485 1.420 14.625 2.500 ;
        RECT  14.395 0.925 14.485 2.500 ;
        RECT  14.240 2.730 14.470 3.455 ;
        RECT  14.255 0.925 14.395 1.650 ;
        RECT  14.205 2.270 14.395 2.500 ;
        RECT  13.295 1.420 14.255 1.650 ;
        RECT  12.955 2.730 14.240 2.960 ;
        RECT  13.795 0.465 14.025 1.190 ;
        RECT  13.635 1.880 13.975 2.415 ;
        RECT  12.900 0.960 13.795 1.190 ;
        RECT  12.320 2.185 13.635 2.415 ;
        RECT  12.955 1.420 13.295 1.835 ;
        RECT  12.725 2.730 12.955 3.250 ;
        RECT  12.670 0.465 12.900 1.190 ;
        RECT  11.755 3.020 12.725 3.250 ;
        RECT  10.350 0.465 12.670 0.695 ;
        RECT  12.090 0.935 12.320 2.705 ;
        RECT  11.525 0.925 11.755 2.585 ;
        RECT  11.310 0.925 11.525 1.155 ;
        RECT  11.295 2.345 11.525 3.210 ;
        RECT  11.035 1.615 11.295 1.955 ;
        RECT  8.945 2.980 11.295 3.210 ;
        RECT  10.805 0.925 11.035 2.750 ;
        RECT  10.670 0.925 10.805 1.265 ;
        RECT  10.515 2.520 10.805 2.750 ;
        RECT  10.420 1.770 10.560 2.110 ;
        RECT  10.190 1.155 10.420 2.110 ;
        RECT  10.120 0.465 10.350 0.925 ;
        RECT  9.405 1.155 10.190 1.385 ;
        RECT  8.555 0.695 10.120 0.925 ;
        RECT  9.175 1.155 9.405 2.750 ;
        RECT  8.865 1.155 9.175 1.385 ;
        RECT  8.715 2.120 8.945 3.210 ;
        RECT  7.335 2.120 8.715 2.350 ;
        RECT  8.325 0.695 8.555 1.860 ;
        RECT  8.255 2.645 8.485 3.455 ;
        RECT  7.565 1.630 8.325 1.860 ;
        RECT  6.630 3.225 8.255 3.455 ;
        RECT  7.825 0.505 8.055 1.315 ;
        RECT  5.095 0.505 7.825 0.735 ;
        RECT  7.105 1.020 7.335 2.985 ;
        RECT  3.575 1.020 7.105 1.250 ;
        RECT  6.290 2.910 6.630 3.455 ;
        RECT  4.730 3.225 6.290 3.455 ;
        RECT  4.390 2.960 4.730 3.455 ;
        RECT  4.020 1.480 4.375 1.770 ;
        RECT  3.115 1.480 4.020 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFKCNQD0BWP7T

MACRO SEDFKCNQD1BWP7T
    CLASS CORE ;
    FOREIGN SEDFKCNQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.570 0.470 18.900 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4581 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.820 6.630 2.100 ;
        RECT  5.380 1.540 5.720 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.765 9.940 2.710 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1782 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 2.370 6.860 2.660 ;
        RECT  4.755 1.485 4.985 2.660 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.085 -0.235 19.040 0.235 ;
        RECT  17.855 -0.235 18.085 1.255 ;
        RECT  16.665 -0.235 17.855 0.235 ;
        RECT  16.325 -0.235 16.665 0.465 ;
        RECT  13.565 -0.235 16.325 0.235 ;
        RECT  13.225 -0.235 13.565 0.730 ;
        RECT  9.845 -0.235 13.225 0.235 ;
        RECT  9.505 -0.235 9.845 0.465 ;
        RECT  4.035 -0.235 9.505 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.085 3.685 19.040 4.155 ;
        RECT  17.855 2.255 18.085 4.155 ;
        RECT  16.680 3.685 17.855 4.155 ;
        RECT  16.340 3.455 16.680 4.155 ;
        RECT  13.720 3.685 16.340 4.155 ;
        RECT  13.360 3.190 13.720 4.155 ;
        RECT  10.025 3.685 13.360 4.155 ;
        RECT  9.685 3.455 10.025 4.155 ;
        RECT  3.940 3.685 9.685 4.155 ;
        RECT  3.580 2.960 3.940 4.155 ;
        RECT  1.290 3.685 3.580 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.620 1.600 18.325 1.940 ;
        RECT  17.390 1.020 17.620 2.795 ;
        RECT  17.385 1.020 17.390 1.250 ;
        RECT  17.385 2.565 17.390 2.795 ;
        RECT  17.155 0.495 17.385 1.250 ;
        RECT  17.155 2.565 17.385 3.380 ;
        RECT  16.930 1.565 17.160 2.310 ;
        RECT  16.635 1.020 17.155 1.250 ;
        RECT  16.765 2.080 16.930 2.310 ;
        RECT  16.535 2.080 16.765 2.995 ;
        RECT  16.405 1.020 16.635 1.830 ;
        RECT  15.210 2.765 16.535 2.995 ;
        RECT  16.120 1.600 16.405 1.830 ;
        RECT  15.810 2.300 16.135 2.530 ;
        RECT  15.810 0.990 16.120 1.220 ;
        RECT  14.470 3.225 15.845 3.455 ;
        RECT  15.580 0.465 15.810 2.530 ;
        RECT  14.025 0.465 15.580 0.695 ;
        RECT  14.980 0.925 15.210 2.995 ;
        RECT  14.485 1.420 14.625 2.500 ;
        RECT  14.395 0.925 14.485 2.500 ;
        RECT  14.240 2.730 14.470 3.455 ;
        RECT  14.255 0.925 14.395 1.650 ;
        RECT  14.205 2.270 14.395 2.500 ;
        RECT  13.295 1.420 14.255 1.650 ;
        RECT  12.955 2.730 14.240 2.960 ;
        RECT  13.795 0.465 14.025 1.190 ;
        RECT  13.635 1.880 13.975 2.415 ;
        RECT  12.900 0.960 13.795 1.190 ;
        RECT  12.320 2.185 13.635 2.415 ;
        RECT  12.955 1.420 13.295 1.835 ;
        RECT  12.725 2.730 12.955 3.250 ;
        RECT  12.670 0.465 12.900 1.190 ;
        RECT  11.755 3.020 12.725 3.250 ;
        RECT  10.350 0.465 12.670 0.695 ;
        RECT  12.090 0.935 12.320 2.705 ;
        RECT  11.525 0.925 11.755 2.585 ;
        RECT  11.310 0.925 11.525 1.155 ;
        RECT  11.295 2.345 11.525 3.210 ;
        RECT  11.035 1.615 11.295 1.955 ;
        RECT  8.945 2.980 11.295 3.210 ;
        RECT  10.805 0.925 11.035 2.750 ;
        RECT  10.670 0.925 10.805 1.265 ;
        RECT  10.515 2.520 10.805 2.750 ;
        RECT  10.420 1.770 10.560 2.110 ;
        RECT  10.190 1.155 10.420 2.110 ;
        RECT  10.120 0.465 10.350 0.925 ;
        RECT  9.405 1.155 10.190 1.385 ;
        RECT  8.555 0.695 10.120 0.925 ;
        RECT  9.175 1.155 9.405 2.750 ;
        RECT  8.865 1.155 9.175 1.385 ;
        RECT  8.715 2.120 8.945 3.210 ;
        RECT  7.335 2.120 8.715 2.350 ;
        RECT  8.325 0.695 8.555 1.860 ;
        RECT  8.255 2.645 8.485 3.455 ;
        RECT  7.565 1.630 8.325 1.860 ;
        RECT  6.630 3.225 8.255 3.455 ;
        RECT  7.825 0.505 8.055 1.315 ;
        RECT  5.095 0.505 7.825 0.735 ;
        RECT  7.105 1.020 7.335 2.985 ;
        RECT  3.575 1.020 7.105 1.250 ;
        RECT  6.290 2.910 6.630 3.455 ;
        RECT  4.730 3.225 6.290 3.455 ;
        RECT  4.390 2.960 4.730 3.455 ;
        RECT  4.020 1.480 4.375 1.770 ;
        RECT  3.115 1.480 4.020 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFKCNQD1BWP7T

MACRO SEDFKCNQD2BWP7T
    CLASS CORE ;
    FOREIGN SEDFKCNQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.645 1.060 18.900 2.730 ;
        RECT  18.620 0.470 18.645 3.310 ;
        RECT  18.415 0.470 18.620 1.290 ;
        RECT  18.415 2.500 18.620 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4581 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2376 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 1.820 6.630 2.100 ;
        RECT  5.380 1.540 5.720 2.100 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.660 1.765 9.940 2.710 ;
        END
    END CP
    PIN CN
        ANTENNAGATEAREA 0.1782 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 2.370 6.860 2.660 ;
        RECT  4.755 1.485 4.985 2.660 ;
        END
    END CN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.365 -0.235 19.600 0.235 ;
        RECT  19.135 -0.235 19.365 1.230 ;
        RECT  17.925 -0.235 19.135 0.235 ;
        RECT  17.695 -0.235 17.925 0.725 ;
        RECT  16.530 -0.235 17.695 0.235 ;
        RECT  16.190 -0.235 16.530 0.465 ;
        RECT  13.565 -0.235 16.190 0.235 ;
        RECT  13.225 -0.235 13.565 0.730 ;
        RECT  9.845 -0.235 13.225 0.235 ;
        RECT  9.505 -0.235 9.845 0.465 ;
        RECT  4.035 -0.235 9.505 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.365 3.685 19.600 4.155 ;
        RECT  19.135 2.250 19.365 4.155 ;
        RECT  17.925 3.685 19.135 4.155 ;
        RECT  17.695 3.195 17.925 4.155 ;
        RECT  16.590 3.685 17.695 4.155 ;
        RECT  16.250 3.455 16.590 4.155 ;
        RECT  13.720 3.685 16.250 4.155 ;
        RECT  13.360 3.190 13.720 4.155 ;
        RECT  10.025 3.685 13.360 4.155 ;
        RECT  9.685 3.455 10.025 4.155 ;
        RECT  3.940 3.685 9.685 4.155 ;
        RECT  3.580 2.960 3.940 4.155 ;
        RECT  1.290 3.685 3.580 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.800 1.600 18.360 1.940 ;
        RECT  17.545 1.020 17.800 2.795 ;
        RECT  16.545 1.020 17.545 1.250 ;
        RECT  17.035 2.565 17.545 2.795 ;
        RECT  16.840 1.565 17.070 2.335 ;
        RECT  16.650 2.105 16.840 2.335 ;
        RECT  16.420 2.105 16.650 2.995 ;
        RECT  16.315 1.020 16.545 1.875 ;
        RECT  15.210 2.765 16.420 2.995 ;
        RECT  16.030 1.645 16.315 1.875 ;
        RECT  15.755 2.300 16.045 2.530 ;
        RECT  15.755 0.990 15.985 1.220 ;
        RECT  15.525 0.465 15.755 2.530 ;
        RECT  14.470 3.225 15.755 3.455 ;
        RECT  14.025 0.465 15.525 0.695 ;
        RECT  14.980 0.925 15.210 2.995 ;
        RECT  14.485 1.420 14.625 2.500 ;
        RECT  14.395 0.925 14.485 2.500 ;
        RECT  14.240 2.730 14.470 3.455 ;
        RECT  14.255 0.925 14.395 1.650 ;
        RECT  14.205 2.270 14.395 2.500 ;
        RECT  13.295 1.420 14.255 1.650 ;
        RECT  12.955 2.730 14.240 2.960 ;
        RECT  13.795 0.465 14.025 1.190 ;
        RECT  13.635 1.880 13.975 2.415 ;
        RECT  12.900 0.960 13.795 1.190 ;
        RECT  12.320 2.185 13.635 2.415 ;
        RECT  12.955 1.420 13.295 1.835 ;
        RECT  12.725 2.730 12.955 3.250 ;
        RECT  12.670 0.465 12.900 1.190 ;
        RECT  11.755 3.020 12.725 3.250 ;
        RECT  10.350 0.465 12.670 0.695 ;
        RECT  12.090 0.935 12.320 2.705 ;
        RECT  11.525 0.925 11.755 2.585 ;
        RECT  11.310 0.925 11.525 1.155 ;
        RECT  11.295 2.345 11.525 3.210 ;
        RECT  11.035 1.615 11.295 1.955 ;
        RECT  8.945 2.980 11.295 3.210 ;
        RECT  10.805 0.925 11.035 2.750 ;
        RECT  10.670 0.925 10.805 1.265 ;
        RECT  10.515 2.520 10.805 2.750 ;
        RECT  10.420 1.770 10.560 2.110 ;
        RECT  10.190 1.155 10.420 2.110 ;
        RECT  10.120 0.465 10.350 0.925 ;
        RECT  9.405 1.155 10.190 1.385 ;
        RECT  8.555 0.695 10.120 0.925 ;
        RECT  9.175 1.155 9.405 2.750 ;
        RECT  8.865 1.155 9.175 1.385 ;
        RECT  8.715 2.120 8.945 3.210 ;
        RECT  7.335 2.120 8.715 2.350 ;
        RECT  8.325 0.695 8.555 1.860 ;
        RECT  8.255 2.645 8.485 3.455 ;
        RECT  7.565 1.630 8.325 1.860 ;
        RECT  6.630 3.225 8.255 3.455 ;
        RECT  7.825 0.505 8.055 1.315 ;
        RECT  5.095 0.505 7.825 0.735 ;
        RECT  7.105 1.020 7.335 2.985 ;
        RECT  3.575 1.020 7.105 1.250 ;
        RECT  6.290 2.910 6.630 3.455 ;
        RECT  4.730 3.225 6.290 3.455 ;
        RECT  4.390 2.960 4.730 3.455 ;
        RECT  4.020 1.480 4.375 1.770 ;
        RECT  3.115 1.480 4.020 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFKCNQD2BWP7T

MACRO SEDFQD0BWP7T
    CLASS CORE ;
    FOREIGN SEDFQD0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.450 0.465 17.780 3.380 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.020 -0.235 17.920 0.235 ;
        RECT  16.680 -0.235 17.020 0.710 ;
        RECT  15.005 -0.235 16.680 0.235 ;
        RECT  14.775 -0.235 15.005 0.520 ;
        RECT  12.445 -0.235 14.775 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.020 3.685 17.920 4.155 ;
        RECT  16.680 3.115 17.020 4.155 ;
        RECT  15.535 3.685 16.680 4.155 ;
        RECT  15.190 3.225 15.535 4.155 ;
        RECT  12.520 3.685 15.190 4.155 ;
        RECT  12.160 3.190 12.520 4.155 ;
        RECT  8.905 3.685 12.160 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.800 1.600 17.205 1.940 ;
        RECT  16.570 1.020 16.800 2.730 ;
        RECT  15.510 1.020 16.570 1.250 ;
        RECT  15.960 2.500 16.570 2.730 ;
        RECT  15.845 1.530 16.075 2.200 ;
        RECT  15.550 1.970 15.845 2.200 ;
        RECT  15.320 1.970 15.550 2.995 ;
        RECT  15.280 1.020 15.510 1.740 ;
        RECT  14.020 2.765 15.320 2.995 ;
        RECT  14.880 1.510 15.280 1.740 ;
        RECT  14.545 0.990 14.980 1.220 ;
        RECT  14.545 2.300 14.840 2.530 ;
        RECT  13.270 3.225 14.570 3.455 ;
        RECT  14.315 0.465 14.545 2.530 ;
        RECT  12.905 0.465 14.315 0.695 ;
        RECT  14.020 0.935 14.085 1.275 ;
        RECT  13.790 0.935 14.020 2.995 ;
        RECT  13.135 0.925 13.365 2.500 ;
        RECT  13.040 2.730 13.270 3.455 ;
        RECT  12.165 1.420 13.135 1.650 ;
        RECT  13.015 2.270 13.135 2.500 ;
        RECT  11.835 2.730 13.040 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.630 1.880 12.835 2.110 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  12.400 1.880 12.630 2.415 ;
        RECT  11.200 2.185 12.400 2.415 ;
        RECT  11.825 1.420 12.165 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFQD0BWP7T

MACRO SEDFQD1BWP7T
    CLASS CORE ;
    FOREIGN SEDFQD1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.450 0.465 17.780 3.295 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 -0.235 17.920 0.235 ;
        RECT  16.735 -0.235 16.965 1.235 ;
        RECT  15.005 -0.235 16.735 0.235 ;
        RECT  14.775 -0.235 15.005 0.520 ;
        RECT  12.445 -0.235 14.775 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 3.685 17.920 4.155 ;
        RECT  16.735 2.255 16.965 4.155 ;
        RECT  15.600 3.685 16.735 4.155 ;
        RECT  15.255 3.225 15.600 4.155 ;
        RECT  12.520 3.685 15.255 4.155 ;
        RECT  12.160 3.190 12.520 4.155 ;
        RECT  8.905 3.685 12.160 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.495 1.600 17.205 1.940 ;
        RECT  16.265 1.020 16.495 2.660 ;
        RECT  16.035 0.495 16.265 1.250 ;
        RECT  16.035 2.430 16.265 3.285 ;
        RECT  15.510 1.020 16.035 1.250 ;
        RECT  15.795 1.530 16.025 2.200 ;
        RECT  15.510 1.970 15.795 2.200 ;
        RECT  15.280 1.020 15.510 1.740 ;
        RECT  15.280 1.970 15.510 2.995 ;
        RECT  14.880 1.510 15.280 1.740 ;
        RECT  14.020 2.765 15.280 2.995 ;
        RECT  14.545 0.990 14.980 1.220 ;
        RECT  14.545 2.300 14.840 2.530 ;
        RECT  13.350 3.225 14.570 3.455 ;
        RECT  14.315 0.465 14.545 2.530 ;
        RECT  12.905 0.465 14.315 0.695 ;
        RECT  14.020 0.935 14.085 1.275 ;
        RECT  13.790 0.935 14.020 2.995 ;
        RECT  13.135 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  12.165 1.420 13.135 1.650 ;
        RECT  13.015 2.270 13.135 2.500 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.630 1.880 12.835 2.110 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  12.400 1.880 12.630 2.415 ;
        RECT  11.200 2.185 12.400 2.415 ;
        RECT  11.825 1.420 12.165 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFQD1BWP7T

MACRO SEDFQD2BWP7T
    CLASS CORE ;
    FOREIGN SEDFQD2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN Q
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.525 1.060 17.780 2.730 ;
        RECT  17.500 0.470 17.525 3.310 ;
        RECT  17.295 0.470 17.500 1.290 ;
        RECT  17.295 2.500 17.500 3.310 ;
        END
    END Q
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 -0.235 18.480 0.235 ;
        RECT  18.015 -0.235 18.245 1.230 ;
        RECT  16.805 -0.235 18.015 0.235 ;
        RECT  16.575 -0.235 16.805 0.725 ;
        RECT  15.410 -0.235 16.575 0.235 ;
        RECT  15.070 -0.235 15.410 0.465 ;
        RECT  12.445 -0.235 15.070 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 3.685 18.480 4.155 ;
        RECT  18.015 2.250 18.245 4.155 ;
        RECT  16.805 3.685 18.015 4.155 ;
        RECT  16.575 3.195 16.805 4.155 ;
        RECT  15.470 3.685 16.575 4.155 ;
        RECT  15.130 3.455 15.470 4.155 ;
        RECT  12.520 3.685 15.130 4.155 ;
        RECT  12.160 3.190 12.520 4.155 ;
        RECT  8.905 3.685 12.160 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.680 1.600 17.240 1.940 ;
        RECT  16.425 1.020 16.680 2.795 ;
        RECT  15.425 1.020 16.425 1.250 ;
        RECT  15.915 2.565 16.425 2.795 ;
        RECT  15.720 1.565 15.950 2.335 ;
        RECT  15.530 2.105 15.720 2.335 ;
        RECT  15.300 2.105 15.530 2.995 ;
        RECT  15.195 1.020 15.425 1.875 ;
        RECT  14.090 2.765 15.300 2.995 ;
        RECT  14.910 1.645 15.195 1.875 ;
        RECT  14.635 2.300 14.925 2.530 ;
        RECT  14.635 0.990 14.865 1.220 ;
        RECT  14.405 0.465 14.635 2.530 ;
        RECT  13.350 3.225 14.635 3.455 ;
        RECT  12.905 0.465 14.405 0.695 ;
        RECT  13.860 0.925 14.090 2.995 ;
        RECT  13.135 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  12.165 1.420 13.135 1.650 ;
        RECT  13.015 2.270 13.135 2.500 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.630 1.880 12.835 2.110 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  12.400 1.880 12.630 2.415 ;
        RECT  11.200 2.185 12.400 2.415 ;
        RECT  11.825 1.420 12.165 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFQD2BWP7T

MACRO SEDFQND0BWP7T
    CLASS CORE ;
    FOREIGN SEDFQND0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.450 0.545 17.780 3.400 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.005 -0.235 17.920 0.235 ;
        RECT  14.775 -0.235 15.005 0.520 ;
        RECT  12.445 -0.235 14.775 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 3.685 17.920 4.155 ;
        RECT  16.735 3.060 16.965 4.155 ;
        RECT  15.560 3.685 16.735 4.155 ;
        RECT  15.215 3.345 15.560 4.155 ;
        RECT  12.520 3.685 15.215 4.155 ;
        RECT  12.160 3.190 12.520 4.155 ;
        RECT  8.905 3.685 12.160 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.935 0.485 17.165 1.940 ;
        RECT  15.605 0.485 16.935 0.715 ;
        RECT  16.320 1.245 16.505 2.730 ;
        RECT  16.275 0.955 16.320 2.730 ;
        RECT  15.980 0.955 16.275 1.475 ;
        RECT  15.980 2.500 16.275 2.730 ;
        RECT  15.815 1.705 16.045 2.200 ;
        RECT  15.555 1.245 15.980 1.475 ;
        RECT  15.510 1.970 15.815 2.200 ;
        RECT  15.375 0.485 15.605 1.005 ;
        RECT  15.325 1.245 15.555 1.740 ;
        RECT  15.280 1.970 15.510 2.995 ;
        RECT  14.980 0.775 15.375 1.005 ;
        RECT  14.880 1.510 15.325 1.740 ;
        RECT  14.085 2.765 15.280 2.995 ;
        RECT  14.545 0.775 14.980 1.220 ;
        RECT  14.545 2.300 14.880 2.530 ;
        RECT  14.315 0.465 14.545 2.530 ;
        RECT  13.350 3.225 14.445 3.455 ;
        RECT  12.905 0.465 14.315 0.695 ;
        RECT  13.835 0.935 14.085 2.995 ;
        RECT  13.135 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  12.165 1.420 13.135 1.650 ;
        RECT  13.015 2.270 13.135 2.500 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.630 1.880 12.835 2.110 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  12.400 1.880 12.630 2.415 ;
        RECT  11.200 2.185 12.400 2.415 ;
        RECT  11.825 1.420 12.165 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFQND0BWP7T

MACRO SEDFQND1BWP7T
    CLASS CORE ;
    FOREIGN SEDFQND1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.920 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.1376 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.450 0.465 17.780 3.295 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.005 -0.235 17.920 0.235 ;
        RECT  14.775 -0.235 15.005 0.520 ;
        RECT  12.445 -0.235 14.775 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.965 3.685 17.920 4.155 ;
        RECT  16.735 2.255 16.965 4.155 ;
        RECT  15.600 3.685 16.735 4.155 ;
        RECT  15.255 3.225 15.600 4.155 ;
        RECT  12.520 3.685 15.255 4.155 ;
        RECT  12.160 3.190 12.520 4.155 ;
        RECT  8.905 3.685 12.160 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.935 0.560 17.165 1.940 ;
        RECT  15.605 0.560 16.935 0.790 ;
        RECT  16.320 1.245 16.505 2.660 ;
        RECT  16.275 1.020 16.320 2.660 ;
        RECT  15.980 1.020 16.275 1.475 ;
        RECT  16.265 2.430 16.275 2.660 ;
        RECT  16.035 2.430 16.265 3.285 ;
        RECT  15.815 1.705 16.045 2.200 ;
        RECT  15.555 1.245 15.980 1.475 ;
        RECT  15.510 1.970 15.815 2.200 ;
        RECT  15.375 0.560 15.605 1.005 ;
        RECT  15.325 1.245 15.555 1.740 ;
        RECT  15.280 1.970 15.510 2.995 ;
        RECT  14.980 0.775 15.375 1.005 ;
        RECT  14.880 1.510 15.325 1.740 ;
        RECT  14.085 2.765 15.280 2.995 ;
        RECT  14.545 0.775 14.980 1.220 ;
        RECT  14.545 2.300 14.880 2.530 ;
        RECT  14.315 0.465 14.545 2.530 ;
        RECT  13.350 3.225 14.445 3.455 ;
        RECT  12.905 0.465 14.315 0.695 ;
        RECT  13.835 0.935 14.085 2.995 ;
        RECT  13.135 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  12.165 1.420 13.135 1.650 ;
        RECT  13.015 2.270 13.135 2.500 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.630 1.880 12.835 2.110 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  12.400 1.880 12.630 2.415 ;
        RECT  11.200 2.185 12.400 2.415 ;
        RECT  11.825 1.420 12.165 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFQND1BWP7T

MACRO SEDFQND2BWP7T
    CLASS CORE ;
    FOREIGN SEDFQND2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.480 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN SI
        ANTENNAGATEAREA 0.1512 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.210 1.540 2.260 ;
        END
    END SI
    PIN SE
        ANTENNAGATEAREA 0.4176 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 2.330 4.340 2.710 ;
        RECT  3.355 1.940 3.695 2.710 ;
        END
    END SE
    PIN QN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.525 1.045 17.780 2.720 ;
        RECT  17.500 0.465 17.525 3.295 ;
        RECT  17.295 0.465 17.500 1.275 ;
        RECT  17.295 2.485 17.500 3.295 ;
        END
    END QN
    PIN E
        ANTENNAGATEAREA 0.4041 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.370 ;
        END
    END E
    PIN D
        ANTENNAGATEAREA 0.2718 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.755 5.460 2.150 ;
        END
    END D
    PIN CP
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.540 1.765 8.820 2.710 ;
        RECT  8.465 1.765 8.540 2.105 ;
        END
    END CP
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 -0.235 18.480 0.235 ;
        RECT  18.015 -0.235 18.245 1.255 ;
        RECT  15.145 -0.235 18.015 0.235 ;
        RECT  14.915 -0.235 15.145 0.520 ;
        RECT  12.445 -0.235 14.915 0.235 ;
        RECT  12.105 -0.235 12.445 0.730 ;
        RECT  8.860 -0.235 12.105 0.235 ;
        RECT  8.520 -0.235 8.860 0.465 ;
        RECT  4.035 -0.235 8.520 0.235 ;
        RECT  3.805 -0.235 4.035 0.785 ;
        RECT  1.250 -0.235 3.805 0.235 ;
        RECT  0.890 -0.235 1.250 0.830 ;
        RECT  0.000 -0.235 0.890 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.245 3.685 18.480 4.155 ;
        RECT  18.015 2.255 18.245 4.155 ;
        RECT  16.805 3.685 18.015 4.155 ;
        RECT  16.575 3.190 16.805 4.155 ;
        RECT  15.600 3.685 16.575 4.155 ;
        RECT  15.255 3.225 15.600 4.155 ;
        RECT  12.520 3.685 15.255 4.155 ;
        RECT  12.160 3.190 12.520 4.155 ;
        RECT  8.905 3.685 12.160 4.155 ;
        RECT  8.565 3.455 8.905 4.155 ;
        RECT  3.985 3.685 8.565 4.155 ;
        RECT  3.625 2.960 3.985 4.155 ;
        RECT  1.290 3.685 3.625 4.155 ;
        RECT  0.930 3.190 1.290 4.155 ;
        RECT  0.000 3.685 0.930 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.775 0.560 17.005 1.940 ;
        RECT  15.605 0.560 16.775 0.790 ;
        RECT  16.275 1.245 16.505 2.660 ;
        RECT  16.270 1.245 16.275 1.475 ;
        RECT  15.970 2.430 16.275 2.660 ;
        RECT  15.930 1.020 16.270 1.475 ;
        RECT  15.815 1.705 16.045 2.200 ;
        RECT  15.555 1.245 15.930 1.475 ;
        RECT  15.510 1.970 15.815 2.200 ;
        RECT  15.375 0.560 15.605 1.005 ;
        RECT  15.325 1.245 15.555 1.740 ;
        RECT  15.280 1.970 15.510 2.995 ;
        RECT  14.860 0.775 15.375 1.005 ;
        RECT  14.860 1.510 15.325 1.740 ;
        RECT  14.085 2.765 15.280 2.995 ;
        RECT  14.590 2.300 14.880 2.530 ;
        RECT  14.590 0.775 14.860 1.220 ;
        RECT  14.360 0.465 14.590 2.530 ;
        RECT  13.350 3.225 14.445 3.455 ;
        RECT  12.905 0.465 14.360 0.695 ;
        RECT  13.835 0.935 14.085 2.995 ;
        RECT  13.135 0.925 13.365 2.500 ;
        RECT  13.120 2.730 13.350 3.455 ;
        RECT  12.165 1.420 13.135 1.650 ;
        RECT  13.015 2.270 13.135 2.500 ;
        RECT  11.835 2.730 13.120 2.960 ;
        RECT  12.675 0.465 12.905 1.190 ;
        RECT  12.630 1.880 12.835 2.110 ;
        RECT  11.780 0.960 12.675 1.190 ;
        RECT  12.400 1.880 12.630 2.415 ;
        RECT  11.200 2.185 12.400 2.415 ;
        RECT  11.825 1.420 12.165 1.835 ;
        RECT  11.605 2.730 11.835 3.250 ;
        RECT  11.550 0.465 11.780 1.190 ;
        RECT  10.540 3.020 11.605 3.250 ;
        RECT  9.320 0.465 11.550 0.695 ;
        RECT  10.970 0.935 11.200 2.650 ;
        RECT  10.765 2.420 10.970 2.650 ;
        RECT  10.310 0.985 10.535 2.625 ;
        RECT  10.305 0.985 10.310 3.210 ;
        RECT  10.190 0.985 10.305 1.220 ;
        RECT  10.080 2.345 10.305 3.210 ;
        RECT  7.775 2.980 10.080 3.210 ;
        RECT  9.825 1.615 10.035 1.955 ;
        RECT  9.595 0.925 9.825 2.670 ;
        RECT  9.550 0.925 9.595 1.265 ;
        RECT  9.320 2.440 9.595 2.670 ;
        RECT  9.300 1.770 9.365 2.110 ;
        RECT  9.090 0.465 9.320 0.925 ;
        RECT  9.070 1.155 9.300 2.110 ;
        RECT  7.735 0.695 9.090 0.925 ;
        RECT  8.235 1.155 9.070 1.385 ;
        RECT  8.235 2.410 8.290 2.750 ;
        RECT  8.005 1.155 8.235 2.750 ;
        RECT  7.545 2.555 7.775 3.210 ;
        RECT  7.505 0.695 7.735 2.165 ;
        RECT  6.180 2.555 7.545 2.785 ;
        RECT  6.640 1.935 7.505 2.165 ;
        RECT  7.085 3.015 7.315 3.360 ;
        RECT  6.945 0.505 7.175 1.315 ;
        RECT  4.800 3.130 7.085 3.360 ;
        RECT  4.540 0.505 6.945 0.735 ;
        RECT  5.950 1.020 6.180 2.785 ;
        RECT  3.575 1.020 5.950 1.250 ;
        RECT  5.725 2.555 5.950 2.785 ;
        RECT  4.570 2.580 4.800 3.360 ;
        RECT  4.025 1.480 4.380 1.770 ;
        RECT  3.115 1.480 4.025 1.710 ;
        RECT  3.345 0.465 3.575 1.250 ;
        RECT  2.415 0.465 3.345 0.695 ;
        RECT  2.885 0.955 3.115 2.890 ;
        RECT  2.695 1.715 2.885 2.055 ;
        RECT  1.850 3.225 2.660 3.455 ;
        RECT  2.185 0.465 2.415 2.930 ;
        RECT  1.620 2.730 1.850 3.455 ;
        RECT  0.465 2.730 1.620 2.960 ;
        RECT  0.235 0.575 0.465 2.960 ;
    END
END SEDFQND2BWP7T

MACRO TAPCELLBWP7T
    CLASS CORE ;
    FOREIGN TAPCELLBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.120 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 -0.235 1.120 0.235 ;
        RECT  0.370 -0.235 0.750 1.140 ;
        RECT  0.000 -0.235 0.370 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 3.685 1.120 4.155 ;
        RECT  0.370 2.610 0.750 4.155 ;
        RECT  0.000 3.685 0.370 4.155 ;
        END
    END VDD
END TAPCELLBWP7T

MACRO TIEHBWP7T
    CLASS CORE ;
    FOREIGN TIEHBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.6850 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.770 1.540 2.710 ;
        RECT  1.260 1.770 1.330 3.425 ;
        RECT  1.090 2.305 1.260 3.425 ;
        END
    END Z
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.400 -0.235 1.680 0.235 ;
        RECT  1.020 -0.235 1.400 1.195 ;
        RECT  0.000 -0.235 1.020 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.680 3.685 1.680 4.155 ;
        RECT  0.300 2.310 0.680 4.155 ;
        RECT  0.000 3.685 0.300 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.370 0.495 0.610 1.955 ;
    END
END TIEHBWP7T

MACRO TIELBWP7T
    CLASS CORE ;
    FOREIGN TIELBWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.680 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.4800 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.000 1.540 2.150 ;
        RECT  1.260 0.495 1.330 2.150 ;
        RECT  1.090 0.495 1.260 1.330 ;
        END
    END ZN
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.680 -0.235 1.680 0.235 ;
        RECT  0.300 -0.235 0.680 1.205 ;
        RECT  0.000 -0.235 0.300 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.400 3.685 1.680 4.155 ;
        RECT  1.020 2.565 1.400 4.155 ;
        RECT  0.000 3.685 1.020 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.370 1.605 0.610 3.400 ;
    END
END TIELBWP7T

MACRO XNR2D0BWP7T
    CLASS CORE ;
    FOREIGN XNR2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.5913 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 0.965 5.460 2.990 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.770 4.340 2.710 ;
        RECT  3.935 1.770 4.060 2.170 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.770 0.980 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.475 -0.235 5.600 0.235 ;
        RECT  5.035 -0.235 5.475 0.465 ;
        RECT  1.365 -0.235 5.035 0.235 ;
        RECT  0.985 -0.235 1.365 0.785 ;
        RECT  0.000 -0.235 0.985 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.680 3.685 5.600 4.155 ;
        RECT  4.300 2.960 4.680 4.155 ;
        RECT  1.320 3.685 4.300 4.155 ;
        RECT  0.940 3.035 1.320 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.640 1.090 4.875 2.140 ;
        RECT  4.455 1.090 4.640 1.360 ;
        RECT  4.215 0.550 4.455 1.360 ;
        RECT  3.215 0.550 4.215 0.785 ;
        RECT  3.675 1.020 3.915 1.255 ;
        RECT  3.690 2.580 3.810 2.920 ;
        RECT  3.675 2.580 3.690 3.420 ;
        RECT  3.445 1.020 3.675 3.420 ;
        RECT  1.845 3.180 3.445 3.420 ;
        RECT  2.975 0.550 3.215 2.870 ;
        RECT  2.695 0.550 2.975 0.785 ;
        RECT  2.795 2.630 2.975 2.870 ;
        RECT  2.505 1.015 2.735 2.370 ;
        RECT  1.825 1.015 2.505 1.255 ;
        RECT  2.325 2.130 2.505 2.370 ;
        RECT  2.085 2.130 2.325 2.920 ;
        RECT  2.025 1.500 2.265 1.900 ;
        RECT  1.515 1.500 2.025 1.740 ;
        RECT  1.645 2.350 1.845 3.420 ;
        RECT  1.605 2.035 1.645 3.420 ;
        RECT  1.305 2.035 1.605 2.580 ;
        RECT  1.245 1.020 1.515 1.740 ;
        RECT  0.380 1.020 1.245 1.255 ;
        RECT  0.380 3.030 0.520 3.270 ;
        RECT  0.140 1.020 0.380 3.270 ;
    END
END XNR2D0BWP7T

MACRO XNR2D1BWP7T
    CLASS CORE ;
    FOREIGN XNR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.040 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1495 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.570 0.465 4.900 3.145 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        RECT  3.420 1.210 3.500 1.850 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.200 0.980 2.150 ;
        RECT  0.580 1.760 0.700 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.130 -0.235 5.040 0.235 ;
        RECT  3.750 -0.235 4.130 0.930 ;
        RECT  1.305 -0.235 3.750 0.235 ;
        RECT  0.925 -0.235 1.305 0.785 ;
        RECT  0.000 -0.235 0.925 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.140 3.685 5.040 4.155 ;
        RECT  3.760 3.245 4.140 4.155 ;
        RECT  1.285 3.685 3.760 4.155 ;
        RECT  0.905 2.890 1.285 4.155 ;
        RECT  0.000 3.685 0.905 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.060 1.620 4.340 3.015 ;
        RECT  2.690 2.785 4.060 3.015 ;
        RECT  3.165 0.545 3.365 0.805 ;
        RECT  3.165 2.325 3.345 2.555 ;
        RECT  2.935 0.545 3.165 2.555 ;
        RECT  1.775 0.545 2.935 0.785 ;
        RECT  2.410 1.015 2.690 3.015 ;
        RECT  2.125 1.015 2.410 1.255 ;
        RECT  2.245 2.695 2.410 3.015 ;
        RECT  1.950 1.555 2.180 2.340 ;
        RECT  1.555 2.110 1.950 2.340 ;
        RECT  1.535 0.545 1.775 1.380 ;
        RECT  1.325 2.110 1.555 2.660 ;
        RECT  1.505 1.150 1.535 1.380 ;
        RECT  1.270 1.150 1.505 1.825 ;
        RECT  0.465 2.420 1.325 2.660 ;
        RECT  0.350 0.630 0.520 0.870 ;
        RECT  0.350 2.420 0.465 2.910 ;
        RECT  0.120 0.630 0.350 2.910 ;
    END
END XNR2D1BWP7T

MACRO XNR2D2BWP7T
    CLASS CORE ;
    FOREIGN XNR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 0.495 6.020 3.325 ;
        RECT  5.480 0.495 5.740 1.305 ;
        RECT  5.530 2.985 5.740 3.325 ;
        END
    END ZN
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.620 1.165 4.900 2.150 ;
        RECT  4.375 1.680 4.620 2.020 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.620 1.540 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 -0.235 6.720 0.235 ;
        RECT  6.250 -0.235 6.490 1.250 ;
        RECT  5.060 -0.235 6.250 0.235 ;
        RECT  4.720 -0.235 5.060 0.670 ;
        RECT  1.185 -0.235 4.720 0.235 ;
        RECT  0.955 -0.235 1.185 0.725 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 3.685 6.720 4.155 ;
        RECT  6.255 2.250 6.490 4.155 ;
        RECT  5.110 3.685 6.255 4.155 ;
        RECT  4.730 3.245 5.110 4.155 ;
        RECT  1.280 3.685 4.730 4.155 ;
        RECT  0.940 3.455 1.280 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.360 1.605 5.475 1.945 ;
        RECT  5.130 1.605 5.360 2.610 ;
        RECT  4.975 2.380 5.130 2.610 ;
        RECT  4.745 2.380 4.975 3.015 ;
        RECT  3.525 2.785 4.745 3.015 ;
        RECT  4.095 2.300 4.355 2.530 ;
        RECT  4.095 1.015 4.300 1.255 ;
        RECT  3.865 0.465 4.095 2.530 ;
        RECT  1.645 0.465 3.865 0.705 ;
        RECT  3.295 0.945 3.525 3.015 ;
        RECT  2.540 0.945 2.820 3.225 ;
        RECT  0.520 2.995 2.540 3.225 ;
        RECT  1.875 0.965 2.175 2.585 ;
        RECT  1.415 0.465 1.645 1.215 ;
        RECT  1.000 0.985 1.415 1.215 ;
        RECT  0.805 0.985 1.000 1.860 ;
        RECT  0.770 0.985 0.805 2.035 ;
        RECT  0.575 1.620 0.770 2.035 ;
        RECT  0.345 2.490 0.520 3.225 ;
        RECT  0.345 0.495 0.465 1.305 ;
        RECT  0.115 0.495 0.345 3.225 ;
    END
END XNR2D2BWP7T

MACRO XNR3D0BWP7T
    CLASS CORE ;
    FOREIGN XNR3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.050 0.465 9.380 2.865 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.210 8.260 2.150 ;
        RECT  7.900 1.210 7.980 1.850 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2502 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        RECT  3.725 1.625 4.060 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.610 -0.235 9.520 0.235 ;
        RECT  8.230 -0.235 8.610 0.790 ;
        RECT  5.720 -0.235 8.230 0.235 ;
        RECT  5.490 -0.235 5.720 0.840 ;
        RECT  4.225 -0.235 5.490 0.235 ;
        RECT  3.845 -0.235 4.225 0.970 ;
        RECT  1.305 -0.235 3.845 0.235 ;
        RECT  0.925 -0.235 1.305 0.975 ;
        RECT  0.000 -0.235 0.925 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.575 3.685 9.520 4.155 ;
        RECT  8.235 3.455 8.575 4.155 ;
        RECT  5.720 3.685 8.235 4.155 ;
        RECT  5.490 3.120 5.720 4.155 ;
        RECT  4.225 3.685 5.490 4.155 ;
        RECT  3.885 3.450 4.225 4.155 ;
        RECT  1.260 3.685 3.885 4.155 ;
        RECT  0.880 2.890 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.570 1.620 8.800 3.070 ;
        RECT  7.130 2.840 8.570 3.070 ;
        RECT  7.645 0.545 7.845 0.805 ;
        RECT  7.645 2.245 7.750 2.585 ;
        RECT  7.415 0.545 7.645 2.585 ;
        RECT  6.265 0.545 7.415 0.785 ;
        RECT  6.900 1.015 7.130 3.070 ;
        RECT  6.615 1.015 6.900 1.255 ;
        RECT  6.705 2.705 6.900 2.935 ;
        RECT  6.440 1.555 6.670 2.340 ;
        RECT  5.530 2.110 6.440 2.340 ;
        RECT  6.025 0.545 6.265 1.380 ;
        RECT  5.995 1.150 6.025 1.380 ;
        RECT  5.760 1.150 5.995 1.825 ;
        RECT  5.300 1.180 5.530 2.890 ;
        RECT  5.240 1.180 5.300 1.410 ;
        RECT  5.260 2.660 5.300 2.890 ;
        RECT  5.030 2.660 5.260 3.405 ;
        RECT  5.010 0.635 5.240 1.410 ;
        RECT  4.660 3.175 5.030 3.405 ;
        RECT  4.660 0.635 5.010 0.865 ;
        RECT  4.800 1.760 4.975 2.100 ;
        RECT  4.570 1.760 4.800 2.945 ;
        RECT  4.295 2.705 4.570 2.945 ;
        RECT  4.055 2.705 4.295 3.220 ;
        RECT  2.845 2.990 4.055 3.220 ;
        RECT  3.085 0.510 3.445 2.760 ;
        RECT  1.835 0.510 3.085 0.740 ;
        RECT  2.605 1.015 2.845 3.220 ;
        RECT  2.325 1.015 2.605 1.255 ;
        RECT  2.285 2.690 2.605 2.930 ;
        RECT  2.140 1.485 2.370 2.420 ;
        RECT  1.880 2.180 2.140 2.420 ;
        RECT  1.650 2.180 1.880 2.620 ;
        RECT  1.605 0.510 1.835 1.775 ;
        RECT  0.470 2.380 1.650 2.620 ;
        RECT  1.390 1.535 1.605 1.775 ;
        RECT  0.230 0.925 0.470 3.165 ;
    END
END XNR3D0BWP7T

MACRO XNR3D1BWP7T
    CLASS CORE ;
    FOREIGN XNR3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.1495 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.050 0.465 9.380 3.145 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.210 8.260 2.150 ;
        RECT  7.900 1.210 7.980 1.850 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4257 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        RECT  3.725 1.625 4.060 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.610 -0.235 9.520 0.235 ;
        RECT  8.230 -0.235 8.610 0.930 ;
        RECT  5.720 -0.235 8.230 0.235 ;
        RECT  5.490 -0.235 5.720 0.840 ;
        RECT  4.225 -0.235 5.490 0.235 ;
        RECT  3.845 -0.235 4.225 0.970 ;
        RECT  1.305 -0.235 3.845 0.235 ;
        RECT  0.925 -0.235 1.305 0.975 ;
        RECT  0.000 -0.235 0.925 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.620 3.685 9.520 4.155 ;
        RECT  8.240 3.245 8.620 4.155 ;
        RECT  5.720 3.685 8.240 4.155 ;
        RECT  5.490 3.120 5.720 4.155 ;
        RECT  4.225 3.685 5.490 4.155 ;
        RECT  3.885 3.450 4.225 4.155 ;
        RECT  1.260 3.685 3.885 4.155 ;
        RECT  0.880 2.890 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.540 1.620 8.820 3.015 ;
        RECT  7.170 2.785 8.540 3.015 ;
        RECT  7.645 0.545 7.845 0.805 ;
        RECT  7.645 2.325 7.825 2.555 ;
        RECT  7.415 0.545 7.645 2.555 ;
        RECT  6.265 0.545 7.415 0.785 ;
        RECT  6.900 1.015 7.170 3.015 ;
        RECT  6.615 1.015 6.900 1.255 ;
        RECT  6.725 2.695 6.900 3.015 ;
        RECT  6.440 1.555 6.670 2.340 ;
        RECT  5.530 2.110 6.440 2.340 ;
        RECT  6.025 0.545 6.265 1.380 ;
        RECT  5.995 1.150 6.025 1.380 ;
        RECT  5.760 1.150 5.995 1.825 ;
        RECT  5.300 1.180 5.530 2.690 ;
        RECT  5.240 1.180 5.300 1.410 ;
        RECT  5.260 2.460 5.300 2.690 ;
        RECT  5.030 2.460 5.260 3.405 ;
        RECT  5.010 0.635 5.240 1.410 ;
        RECT  4.660 3.175 5.030 3.405 ;
        RECT  4.660 0.635 5.010 0.865 ;
        RECT  4.800 1.760 4.975 2.100 ;
        RECT  4.570 1.760 4.800 2.735 ;
        RECT  4.295 2.495 4.570 2.735 ;
        RECT  4.055 2.495 4.295 3.220 ;
        RECT  2.845 2.980 4.055 3.220 ;
        RECT  3.085 0.510 3.445 2.745 ;
        RECT  1.835 0.510 3.085 0.740 ;
        RECT  2.605 1.015 2.845 3.220 ;
        RECT  2.325 1.015 2.605 1.255 ;
        RECT  2.285 2.690 2.605 2.930 ;
        RECT  2.140 1.600 2.370 2.420 ;
        RECT  1.880 2.180 2.140 2.420 ;
        RECT  1.650 2.180 1.880 2.620 ;
        RECT  1.605 0.510 1.835 1.905 ;
        RECT  0.470 2.380 1.650 2.620 ;
        RECT  1.390 1.665 1.605 1.905 ;
        RECT  0.230 0.925 0.470 3.165 ;
    END
END XNR3D1BWP7T

MACRO XNR3D2BWP7T
    CLASS CORE ;
    FOREIGN XNR3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.130 0.705 9.380 2.635 ;
        RECT  9.100 0.480 9.130 3.375 ;
        RECT  8.890 0.480 9.100 0.935 ;
        RECT  8.890 2.405 9.100 3.375 ;
        END
    END ZN
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.680 8.260 2.710 ;
        RECT  7.635 1.680 7.980 2.020 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.595 1.210 1.030 2.100 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.850 -0.235 10.080 0.235 ;
        RECT  9.610 -0.235 9.850 1.225 ;
        RECT  8.405 -0.235 9.610 0.235 ;
        RECT  8.175 -0.235 8.405 0.725 ;
        RECT  5.335 -0.235 8.175 0.235 ;
        RECT  5.105 -0.235 5.335 1.085 ;
        RECT  3.970 -0.235 5.105 0.235 ;
        RECT  3.550 -0.235 3.970 0.670 ;
        RECT  1.260 -0.235 3.550 0.235 ;
        RECT  0.880 -0.235 1.260 0.830 ;
        RECT  0.000 -0.235 0.880 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.850 3.685 10.080 4.155 ;
        RECT  9.610 2.510 9.850 4.155 ;
        RECT  8.310 3.685 9.610 4.155 ;
        RECT  7.930 2.960 8.310 4.155 ;
        RECT  5.375 3.685 7.930 4.155 ;
        RECT  5.145 2.760 5.375 4.155 ;
        RECT  4.080 3.685 5.145 4.155 ;
        RECT  3.740 3.450 4.080 4.155 ;
        RECT  1.280 3.685 3.740 4.155 ;
        RECT  0.940 3.250 1.280 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.550 1.210 8.830 2.080 ;
        RECT  7.945 1.210 8.550 1.440 ;
        RECT  7.715 0.465 7.945 1.440 ;
        RECT  6.810 0.465 7.715 0.695 ;
        RECT  7.405 2.400 7.510 2.740 ;
        RECT  7.405 0.965 7.485 1.305 ;
        RECT  7.355 0.965 7.405 2.740 ;
        RECT  7.125 0.965 7.355 3.455 ;
        RECT  5.835 3.225 7.125 3.455 ;
        RECT  6.535 0.465 6.810 2.830 ;
        RECT  6.470 2.585 6.535 2.830 ;
        RECT  6.055 1.315 6.285 1.870 ;
        RECT  4.615 1.315 6.055 1.545 ;
        RECT  5.625 2.210 5.835 3.455 ;
        RECT  5.605 1.775 5.625 3.455 ;
        RECT  5.395 1.775 5.605 2.440 ;
        RECT  5.230 1.775 5.395 2.010 ;
        RECT  4.520 2.990 4.860 3.455 ;
        RECT  4.385 0.875 4.615 2.585 ;
        RECT  3.755 2.990 4.520 3.220 ;
        RECT  3.525 2.760 3.755 3.220 ;
        RECT  2.625 2.760 3.525 2.990 ;
        RECT  3.210 2.300 3.320 2.530 ;
        RECT  3.135 0.790 3.210 2.530 ;
        RECT  2.980 0.465 3.135 2.530 ;
        RECT  2.905 0.465 2.980 1.155 ;
        RECT  1.755 0.465 2.905 0.695 ;
        RECT  2.395 0.935 2.625 2.990 ;
        RECT  2.120 0.935 2.395 1.175 ;
        RECT  2.260 2.430 2.395 2.660 ;
        RECT  1.840 3.225 2.370 3.455 ;
        RECT  2.030 1.485 2.165 1.830 ;
        RECT  1.935 1.485 2.030 2.560 ;
        RECT  1.800 1.600 1.935 2.560 ;
        RECT  1.610 2.790 1.840 3.455 ;
        RECT  0.365 2.330 1.800 2.560 ;
        RECT  1.525 0.465 1.755 1.320 ;
        RECT  0.685 2.790 1.610 3.020 ;
        RECT  1.495 1.090 1.525 1.320 ;
        RECT  1.265 1.090 1.495 1.825 ;
        RECT  0.455 2.790 0.685 3.380 ;
        RECT  0.365 0.585 0.520 0.830 ;
        RECT  0.135 0.585 0.365 2.560 ;
    END
END XNR3D2BWP7T

MACRO XNR4D0BWP7T
    CLASS CORE ;
    FOREIGN XNR4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 0.765 8.260 2.535 ;
        RECT  7.880 0.765 7.980 0.995 ;
        RECT  7.880 2.295 7.980 2.535 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.210 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.170 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 1.600 9.205 1.960 ;
        RECT  8.540 1.210 8.820 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.210 12.180 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 -0.235 12.880 0.235 ;
        RECT  11.695 -0.235 11.930 0.980 ;
        RECT  9.040 -0.235 11.695 0.235 ;
        RECT  8.660 -0.235 9.040 0.970 ;
        RECT  5.545 -0.235 8.660 0.235 ;
        RECT  5.315 -0.235 5.545 1.165 ;
        RECT  4.190 -0.235 5.315 0.235 ;
        RECT  3.810 -0.235 4.190 0.825 ;
        RECT  1.295 -0.235 3.810 0.235 ;
        RECT  0.915 -0.235 1.295 0.830 ;
        RECT  0.000 -0.235 0.915 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 3.685 12.880 4.155 ;
        RECT  11.695 3.025 11.930 4.155 ;
        RECT  8.980 3.685 11.695 4.155 ;
        RECT  8.615 3.445 8.980 4.155 ;
        RECT  5.620 3.685 8.615 4.155 ;
        RECT  5.240 2.565 5.620 4.155 ;
        RECT  4.125 3.685 5.240 4.155 ;
        RECT  3.895 3.195 4.125 4.155 ;
        RECT  1.250 3.685 3.895 4.155 ;
        RECT  0.870 3.060 1.250 4.155 ;
        RECT  0.000 3.685 0.870 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.410 0.670 12.650 3.230 ;
        RECT  11.500 2.510 12.410 2.750 ;
        RECT  11.270 2.035 11.500 2.750 ;
        RECT  11.235 0.465 11.465 1.755 ;
        RECT  10.690 2.035 11.270 2.275 ;
        RECT  9.770 0.465 11.235 0.695 ;
        RECT  10.460 1.820 10.690 2.275 ;
        RECT  10.230 0.945 10.505 1.185 ;
        RECT  10.230 2.585 10.505 2.815 ;
        RECT  10.000 0.945 10.230 2.995 ;
        RECT  7.470 2.765 10.000 2.995 ;
        RECT  9.540 0.465 9.770 2.530 ;
        RECT  9.400 0.725 9.540 0.955 ;
        RECT  9.405 2.300 9.540 2.530 ;
        RECT  7.000 3.225 7.850 3.455 ;
        RECT  7.230 0.465 7.470 2.995 ;
        RECT  6.005 0.465 7.230 0.695 ;
        RECT  6.770 0.945 7.000 3.455 ;
        RECT  6.445 0.945 6.770 1.185 ;
        RECT  6.460 2.610 6.770 2.840 ;
        RECT  6.275 1.775 6.505 2.195 ;
        RECT  4.945 1.965 6.275 2.195 ;
        RECT  5.775 0.465 6.005 1.725 ;
        RECT  5.480 1.475 5.775 1.725 ;
        RECT  4.705 0.910 4.945 2.695 ;
        RECT  4.540 0.910 4.705 1.140 ;
        RECT  4.540 2.465 4.705 2.695 ;
        RECT  4.250 1.600 4.425 1.940 ;
        RECT  4.020 1.600 4.250 2.675 ;
        RECT  3.710 2.445 4.020 2.675 ;
        RECT  3.480 2.445 3.710 3.045 ;
        RECT  2.775 2.815 3.480 3.045 ;
        RECT  3.020 0.465 3.250 2.585 ;
        RECT  1.755 0.465 3.020 0.695 ;
        RECT  2.545 0.975 2.775 3.045 ;
        RECT  2.205 0.975 2.545 1.215 ;
        RECT  2.205 2.555 2.545 2.785 ;
        RECT  2.020 1.855 2.250 2.275 ;
        RECT  1.530 2.045 2.020 2.275 ;
        RECT  1.530 0.465 1.755 1.290 ;
        RECT  1.525 0.465 1.530 1.815 ;
        RECT  1.300 2.045 1.530 2.610 ;
        RECT  1.300 1.060 1.525 1.815 ;
        RECT  0.520 2.380 1.300 2.610 ;
        RECT  0.375 0.585 0.520 0.830 ;
        RECT  0.375 2.380 0.520 3.060 ;
        RECT  0.135 0.585 0.375 3.060 ;
    END
END XNR4D0BWP7T

MACRO XNR4D1BWP7T
    CLASS CORE ;
    FOREIGN XNR4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.0360 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 0.765 8.260 2.535 ;
        RECT  7.880 0.765 7.980 0.995 ;
        RECT  7.880 2.295 7.980 2.535 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.210 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.170 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 1.600 9.205 1.960 ;
        RECT  8.540 1.210 8.820 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.210 12.180 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 -0.235 12.880 0.235 ;
        RECT  11.695 -0.235 11.930 0.980 ;
        RECT  9.040 -0.235 11.695 0.235 ;
        RECT  8.660 -0.235 9.040 0.970 ;
        RECT  5.545 -0.235 8.660 0.235 ;
        RECT  5.315 -0.235 5.545 1.165 ;
        RECT  4.190 -0.235 5.315 0.235 ;
        RECT  3.810 -0.235 4.190 0.825 ;
        RECT  1.295 -0.235 3.810 0.235 ;
        RECT  0.915 -0.235 1.295 0.830 ;
        RECT  0.000 -0.235 0.915 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 3.685 12.880 4.155 ;
        RECT  11.695 3.025 11.930 4.155 ;
        RECT  8.980 3.685 11.695 4.155 ;
        RECT  8.615 3.445 8.980 4.155 ;
        RECT  5.620 3.685 8.615 4.155 ;
        RECT  5.240 2.565 5.620 4.155 ;
        RECT  4.125 3.685 5.240 4.155 ;
        RECT  3.895 3.195 4.125 4.155 ;
        RECT  1.250 3.685 3.895 4.155 ;
        RECT  0.870 3.060 1.250 4.155 ;
        RECT  0.000 3.685 0.870 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.410 0.670 12.650 3.230 ;
        RECT  11.500 2.510 12.410 2.750 ;
        RECT  11.270 2.035 11.500 2.750 ;
        RECT  11.235 0.465 11.465 1.755 ;
        RECT  10.690 2.035 11.270 2.275 ;
        RECT  9.770 0.465 11.235 0.695 ;
        RECT  10.460 1.820 10.690 2.275 ;
        RECT  10.230 0.945 10.505 1.185 ;
        RECT  10.230 2.585 10.505 2.815 ;
        RECT  10.000 0.945 10.230 2.995 ;
        RECT  7.470 2.765 10.000 2.995 ;
        RECT  9.540 0.465 9.770 2.530 ;
        RECT  9.400 0.725 9.540 0.955 ;
        RECT  9.405 2.300 9.540 2.530 ;
        RECT  7.000 3.225 7.850 3.455 ;
        RECT  7.230 0.465 7.470 2.995 ;
        RECT  6.005 0.465 7.230 0.695 ;
        RECT  6.770 0.945 7.000 3.455 ;
        RECT  6.445 0.945 6.770 1.185 ;
        RECT  6.460 2.610 6.770 2.840 ;
        RECT  6.275 1.775 6.505 2.195 ;
        RECT  4.945 1.965 6.275 2.195 ;
        RECT  5.775 0.465 6.005 1.725 ;
        RECT  5.480 1.475 5.775 1.725 ;
        RECT  4.705 0.910 4.945 2.695 ;
        RECT  4.540 0.910 4.705 1.140 ;
        RECT  4.540 2.465 4.705 2.695 ;
        RECT  4.250 1.600 4.425 1.940 ;
        RECT  4.020 1.600 4.250 2.675 ;
        RECT  3.710 2.445 4.020 2.675 ;
        RECT  3.480 2.445 3.710 3.045 ;
        RECT  2.775 2.815 3.480 3.045 ;
        RECT  3.020 0.465 3.250 2.585 ;
        RECT  1.755 0.465 3.020 0.695 ;
        RECT  2.545 0.985 2.775 3.045 ;
        RECT  2.205 0.985 2.545 1.225 ;
        RECT  2.205 2.555 2.545 2.785 ;
        RECT  2.020 1.865 2.250 2.285 ;
        RECT  1.530 2.055 2.020 2.285 ;
        RECT  1.530 0.465 1.755 1.290 ;
        RECT  1.525 0.465 1.530 1.825 ;
        RECT  1.300 2.055 1.530 2.610 ;
        RECT  1.300 1.060 1.525 1.825 ;
        RECT  0.520 2.380 1.300 2.610 ;
        RECT  0.375 0.585 0.520 0.830 ;
        RECT  0.375 2.380 0.520 3.060 ;
        RECT  0.135 0.585 0.375 3.060 ;
    END
END XNR4D1BWP7T

MACRO XNR4D2BWP7T
    CLASS CORE ;
    FOREIGN XNR4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN ZN
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 0.765 8.940 0.995 ;
        RECT  8.820 2.295 8.940 2.530 ;
        RECT  8.540 0.765 8.820 2.530 ;
        END
    END ZN
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.210 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.780 2.170 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.655 1.210 9.940 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.460 1.210 12.740 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.490 -0.235 13.440 0.235 ;
        RECT  12.255 -0.235 12.490 0.980 ;
        RECT  9.700 -0.235 12.255 0.235 ;
        RECT  9.320 -0.235 9.700 0.970 ;
        RECT  8.220 -0.235 9.320 0.235 ;
        RECT  7.880 -0.235 8.220 0.725 ;
        RECT  5.545 -0.235 7.880 0.235 ;
        RECT  5.315 -0.235 5.545 1.165 ;
        RECT  4.190 -0.235 5.315 0.235 ;
        RECT  3.810 -0.235 4.190 0.825 ;
        RECT  1.295 -0.235 3.810 0.235 ;
        RECT  0.915 -0.235 1.295 0.830 ;
        RECT  0.000 -0.235 0.915 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.490 3.685 13.440 4.155 ;
        RECT  12.255 3.025 12.490 4.155 ;
        RECT  9.700 3.685 12.255 4.155 ;
        RECT  9.335 3.250 9.700 4.155 ;
        RECT  8.220 3.685 9.335 4.155 ;
        RECT  7.880 3.250 8.220 4.155 ;
        RECT  5.620 3.685 7.880 4.155 ;
        RECT  5.240 2.565 5.620 4.155 ;
        RECT  4.125 3.685 5.240 4.155 ;
        RECT  3.895 3.195 4.125 4.155 ;
        RECT  1.250 3.685 3.895 4.155 ;
        RECT  0.870 3.060 1.250 4.155 ;
        RECT  0.000 3.685 0.870 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.970 0.670 13.210 3.230 ;
        RECT  12.060 2.510 12.970 2.750 ;
        RECT  11.830 2.035 12.060 2.750 ;
        RECT  12.025 1.195 12.055 1.755 ;
        RECT  11.825 0.465 12.025 1.755 ;
        RECT  11.385 2.035 11.830 2.275 ;
        RECT  11.795 0.465 11.825 1.425 ;
        RECT  10.465 0.465 11.795 0.695 ;
        RECT  11.155 1.820 11.385 2.275 ;
        RECT  10.925 0.945 11.200 1.185 ;
        RECT  10.925 2.585 11.200 2.815 ;
        RECT  10.695 0.945 10.925 3.020 ;
        RECT  8.140 2.790 10.695 3.020 ;
        RECT  10.235 0.465 10.465 2.560 ;
        RECT  10.095 0.725 10.235 0.955 ;
        RECT  10.100 2.330 10.235 2.560 ;
        RECT  7.900 1.090 8.140 3.020 ;
        RECT  7.470 1.090 7.900 1.330 ;
        RECT  7.235 2.430 7.900 2.770 ;
        RECT  7.000 1.600 7.655 1.940 ;
        RECT  7.230 0.465 7.470 1.330 ;
        RECT  6.005 0.465 7.230 0.695 ;
        RECT  6.770 0.945 7.000 2.840 ;
        RECT  6.445 0.945 6.770 1.185 ;
        RECT  6.460 2.610 6.770 2.840 ;
        RECT  6.275 1.775 6.505 2.195 ;
        RECT  4.945 1.965 6.275 2.195 ;
        RECT  5.775 0.465 6.005 1.725 ;
        RECT  5.480 1.475 5.775 1.725 ;
        RECT  4.705 0.910 4.945 2.695 ;
        RECT  4.540 0.910 4.705 1.140 ;
        RECT  4.540 2.465 4.705 2.695 ;
        RECT  4.250 1.600 4.425 1.940 ;
        RECT  4.020 1.600 4.250 2.675 ;
        RECT  3.710 2.445 4.020 2.675 ;
        RECT  3.480 2.445 3.710 3.045 ;
        RECT  2.775 2.815 3.480 3.045 ;
        RECT  3.020 0.465 3.250 2.585 ;
        RECT  1.755 0.465 3.020 0.695 ;
        RECT  2.545 0.975 2.775 3.045 ;
        RECT  2.205 0.975 2.545 1.215 ;
        RECT  2.205 2.555 2.545 2.785 ;
        RECT  2.020 1.865 2.250 2.285 ;
        RECT  1.530 2.055 2.020 2.285 ;
        RECT  1.530 0.465 1.755 1.290 ;
        RECT  1.525 0.465 1.530 1.825 ;
        RECT  1.300 2.055 1.530 2.610 ;
        RECT  1.300 1.060 1.525 1.825 ;
        RECT  0.520 2.380 1.300 2.610 ;
        RECT  0.375 0.585 0.520 0.830 ;
        RECT  0.375 2.380 0.520 3.060 ;
        RECT  0.135 0.585 0.375 3.060 ;
    END
END XNR4D2BWP7T

MACRO XOR2D0BWP7T
    CLASS CORE ;
    FOREIGN XOR2D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.6016 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 0.965 5.460 3.200 ;
        RECT  5.130 0.965 5.180 1.305 ;
        RECT  5.065 2.960 5.180 3.200 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.770 4.340 2.710 ;
        RECT  3.970 1.770 4.060 2.220 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.660 1.770 0.700 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.460 -0.235 5.600 0.235 ;
        RECT  4.980 -0.235 5.460 0.475 ;
        RECT  1.335 -0.235 4.980 0.235 ;
        RECT  0.955 -0.235 1.335 0.950 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.675 3.685 5.600 4.155 ;
        RECT  4.295 3.005 4.675 4.155 ;
        RECT  1.330 3.685 4.295 4.155 ;
        RECT  0.950 2.975 1.330 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.885 1.960 4.925 2.300 ;
        RECT  4.655 1.145 4.885 2.300 ;
        RECT  4.235 1.145 4.655 1.385 ;
        RECT  3.995 0.465 4.235 1.385 ;
        RECT  3.265 0.465 3.995 0.705 ;
        RECT  3.735 2.940 3.875 3.455 ;
        RECT  3.495 0.965 3.735 3.455 ;
        RECT  1.800 3.215 3.495 3.455 ;
        RECT  3.035 0.465 3.265 2.870 ;
        RECT  2.605 0.465 3.035 0.705 ;
        RECT  2.765 2.630 3.035 2.870 ;
        RECT  2.555 0.950 2.795 2.400 ;
        RECT  2.130 0.950 2.555 1.180 ;
        RECT  2.290 2.170 2.555 2.400 ;
        RECT  2.050 2.170 2.290 2.920 ;
        RECT  2.020 1.455 2.255 1.940 ;
        RECT  1.890 0.560 2.130 1.180 ;
        RECT  1.560 1.960 1.565 3.455 ;
        RECT  1.335 1.960 1.560 2.640 ;
        RECT  1.220 1.250 1.460 1.685 ;
        RECT  0.470 1.250 1.220 1.490 ;
        RECT  0.370 0.965 0.470 1.490 ;
        RECT  0.370 2.615 0.470 2.955 ;
        RECT  0.140 0.965 0.370 2.955 ;
        RECT  1.460 1.455 2.020 1.685 ;
        RECT  1.565 2.405 1.800 3.455 ;
    END
END XOR2D0BWP7T

MACRO XOR2D1BWP7T
    CLASS CORE ;
    FOREIGN XOR2D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.600 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1582 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.180 0.470 5.460 3.090 ;
        RECT  5.130 0.470 5.180 1.285 ;
        RECT  5.120 2.245 5.180 3.090 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.570 4.340 2.710 ;
        RECT  3.970 1.570 4.060 1.910 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4599 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.770 0.980 2.710 ;
        RECT  0.660 1.770 0.700 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.795 -0.235 5.600 0.235 ;
        RECT  4.415 -0.235 4.795 0.750 ;
        RECT  1.335 -0.235 4.415 0.235 ;
        RECT  0.955 -0.235 1.335 0.985 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.675 3.685 5.600 4.155 ;
        RECT  4.295 3.005 4.675 4.155 ;
        RECT  1.330 3.685 4.295 4.155 ;
        RECT  0.950 2.975 1.330 4.155 ;
        RECT  0.000 3.685 0.950 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.885 1.610 4.925 1.950 ;
        RECT  4.655 1.040 4.885 1.950 ;
        RECT  4.185 1.040 4.655 1.270 ;
        RECT  3.955 0.465 4.185 1.270 ;
        RECT  3.255 0.465 3.955 0.695 ;
        RECT  3.725 2.940 3.845 3.455 ;
        RECT  3.485 0.965 3.725 3.455 ;
        RECT  1.800 3.215 3.485 3.455 ;
        RECT  3.025 0.465 3.255 2.870 ;
        RECT  2.605 0.465 3.025 0.695 ;
        RECT  2.765 2.630 3.025 2.870 ;
        RECT  2.555 0.950 2.795 2.400 ;
        RECT  2.130 0.950 2.555 1.180 ;
        RECT  2.290 2.170 2.555 2.400 ;
        RECT  2.050 2.170 2.290 2.920 ;
        RECT  2.020 1.455 2.255 1.940 ;
        RECT  1.890 0.560 2.130 1.180 ;
        RECT  1.560 1.960 1.565 3.455 ;
        RECT  1.335 1.960 1.560 2.640 ;
        RECT  1.220 1.250 1.460 1.685 ;
        RECT  0.470 1.250 1.220 1.490 ;
        RECT  0.370 0.835 0.470 1.490 ;
        RECT  0.370 2.580 0.470 2.920 ;
        RECT  0.140 0.835 0.370 2.920 ;
        RECT  1.460 1.455 2.020 1.685 ;
        RECT  1.565 2.405 1.800 3.455 ;
    END
END XOR2D1BWP7T

MACRO XOR2D2BWP7T
    CLASS CORE ;
    FOREIGN XOR2D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.720 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.740 1.140 6.020 3.040 ;
        RECT  5.500 0.480 5.740 1.400 ;
        RECT  5.500 2.800 5.740 3.365 ;
        END
    END Z
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.590 1.210 4.900 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4905 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.260 1.630 1.540 2.710 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 -0.235 6.720 0.235 ;
        RECT  6.250 -0.235 6.490 1.290 ;
        RECT  5.095 -0.235 6.250 0.235 ;
        RECT  4.715 -0.235 5.095 0.675 ;
        RECT  1.185 -0.235 4.715 0.235 ;
        RECT  0.955 -0.235 1.185 0.725 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 3.685 6.720 4.155 ;
        RECT  6.250 2.255 6.490 4.155 ;
        RECT  5.085 3.685 6.250 4.155 ;
        RECT  4.705 3.250 5.085 4.155 ;
        RECT  1.280 3.685 4.705 4.155 ;
        RECT  0.940 3.455 1.280 4.155 ;
        RECT  0.000 3.685 0.940 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.365 1.630 5.495 1.970 ;
        RECT  5.135 1.630 5.365 2.610 ;
        RECT  4.995 2.380 5.135 2.610 ;
        RECT  4.765 2.380 4.995 3.010 ;
        RECT  3.590 2.780 4.765 3.010 ;
        RECT  4.010 0.465 4.350 2.530 ;
        RECT  1.645 0.465 4.010 0.695 ;
        RECT  3.295 0.965 3.590 3.010 ;
        RECT  2.570 0.965 2.810 3.330 ;
        RECT  1.915 3.090 2.570 3.330 ;
        RECT  1.875 0.965 2.180 2.625 ;
        RECT  1.685 2.985 1.915 3.330 ;
        RECT  0.470 2.985 1.685 3.225 ;
        RECT  1.415 0.465 1.645 1.210 ;
        RECT  0.985 0.980 1.415 1.210 ;
        RECT  0.755 0.980 0.985 2.020 ;
        RECT  0.605 1.680 0.755 2.020 ;
        RECT  0.370 2.330 0.470 3.440 ;
        RECT  0.370 0.495 0.465 1.305 ;
        RECT  0.140 0.495 0.370 3.440 ;
    END
END XOR2D2BWP7T

MACRO XOR3D0BWP7T
    CLASS CORE ;
    FOREIGN XOR3D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5747 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.050 0.465 9.380 2.970 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.210 8.260 2.150 ;
        RECT  7.900 1.210 7.980 1.850 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        RECT  3.740 1.655 4.060 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.610 -0.235 9.520 0.235 ;
        RECT  8.230 -0.235 8.610 0.860 ;
        RECT  5.720 -0.235 8.230 0.235 ;
        RECT  5.490 -0.235 5.720 0.840 ;
        RECT  4.230 -0.235 5.490 0.235 ;
        RECT  3.850 -0.235 4.230 0.830 ;
        RECT  1.285 -0.235 3.850 0.235 ;
        RECT  0.905 -0.235 1.285 0.830 ;
        RECT  0.000 -0.235 0.905 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.575 3.685 9.520 4.155 ;
        RECT  8.235 3.245 8.575 4.155 ;
        RECT  5.720 3.685 8.235 4.155 ;
        RECT  5.490 3.120 5.720 4.155 ;
        RECT  4.225 3.685 5.490 4.155 ;
        RECT  3.865 3.450 4.225 4.155 ;
        RECT  1.260 3.685 3.865 4.155 ;
        RECT  0.880 3.155 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.540 1.620 8.820 3.015 ;
        RECT  7.170 2.785 8.540 3.015 ;
        RECT  7.645 0.545 7.845 0.805 ;
        RECT  7.645 2.325 7.815 2.555 ;
        RECT  7.415 0.545 7.645 2.555 ;
        RECT  6.265 0.545 7.415 0.785 ;
        RECT  6.900 1.015 7.170 3.015 ;
        RECT  6.615 1.015 6.900 1.255 ;
        RECT  6.725 2.550 6.900 2.780 ;
        RECT  6.440 1.555 6.670 2.285 ;
        RECT  5.530 2.055 6.440 2.285 ;
        RECT  6.025 0.545 6.265 1.380 ;
        RECT  5.995 1.150 6.025 1.380 ;
        RECT  5.760 1.150 5.995 1.825 ;
        RECT  5.300 1.180 5.530 2.690 ;
        RECT  5.240 1.180 5.300 1.410 ;
        RECT  5.260 2.460 5.300 2.690 ;
        RECT  5.030 2.460 5.260 3.405 ;
        RECT  5.010 0.635 5.240 1.410 ;
        RECT  4.660 3.175 5.030 3.405 ;
        RECT  4.660 0.635 5.010 0.865 ;
        RECT  4.800 1.760 4.975 2.100 ;
        RECT  4.570 1.760 4.800 2.735 ;
        RECT  4.295 2.495 4.570 2.735 ;
        RECT  4.065 2.495 4.295 3.220 ;
        RECT  2.825 2.990 4.065 3.220 ;
        RECT  3.195 0.520 3.445 2.755 ;
        RECT  1.845 0.520 3.195 0.760 ;
        RECT  3.105 2.525 3.195 2.755 ;
        RECT  2.585 1.000 2.825 3.220 ;
        RECT  2.345 1.000 2.585 1.240 ;
        RECT  2.345 2.670 2.585 2.910 ;
        RECT  2.075 1.680 2.315 2.360 ;
        RECT  1.845 2.130 2.075 2.775 ;
        RECT  1.625 0.520 1.845 1.415 ;
        RECT  0.470 2.545 1.845 2.775 ;
        RECT  1.605 0.520 1.625 1.980 ;
        RECT  1.385 1.175 1.605 1.980 ;
        RECT  0.380 0.560 0.480 0.900 ;
        RECT  0.380 2.545 0.470 3.440 ;
        RECT  0.140 0.560 0.380 3.440 ;
    END
END XOR3D0BWP7T

MACRO XOR3D1BWP7T
    CLASS CORE ;
    FOREIGN XOR3D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.520 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.1495 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.050 0.465 9.380 3.145 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.210 8.260 2.150 ;
        RECT  7.900 1.210 7.980 1.850 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.060 1.210 4.340 2.150 ;
        RECT  3.740 1.655 4.060 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.610 -0.235 9.520 0.235 ;
        RECT  8.230 -0.235 8.610 0.930 ;
        RECT  5.720 -0.235 8.230 0.235 ;
        RECT  5.490 -0.235 5.720 0.840 ;
        RECT  4.230 -0.235 5.490 0.235 ;
        RECT  3.850 -0.235 4.230 0.830 ;
        RECT  1.285 -0.235 3.850 0.235 ;
        RECT  0.905 -0.235 1.285 0.830 ;
        RECT  0.000 -0.235 0.905 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.620 3.685 9.520 4.155 ;
        RECT  8.240 3.245 8.620 4.155 ;
        RECT  5.720 3.685 8.240 4.155 ;
        RECT  5.490 3.120 5.720 4.155 ;
        RECT  4.225 3.685 5.490 4.155 ;
        RECT  3.865 3.450 4.225 4.155 ;
        RECT  1.260 3.685 3.865 4.155 ;
        RECT  0.880 3.155 1.260 4.155 ;
        RECT  0.000 3.685 0.880 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.540 1.620 8.820 3.015 ;
        RECT  7.170 2.785 8.540 3.015 ;
        RECT  7.645 0.545 7.845 0.805 ;
        RECT  7.645 2.325 7.825 2.555 ;
        RECT  7.415 0.545 7.645 2.555 ;
        RECT  6.265 0.545 7.415 0.785 ;
        RECT  6.900 1.015 7.170 3.015 ;
        RECT  6.615 1.015 6.900 1.255 ;
        RECT  6.725 2.695 6.900 3.015 ;
        RECT  6.440 1.555 6.670 2.340 ;
        RECT  5.530 2.110 6.440 2.340 ;
        RECT  6.025 0.545 6.265 1.380 ;
        RECT  5.995 1.150 6.025 1.380 ;
        RECT  5.760 1.150 5.995 1.825 ;
        RECT  5.300 1.180 5.530 2.690 ;
        RECT  5.240 1.180 5.300 1.410 ;
        RECT  5.260 2.460 5.300 2.690 ;
        RECT  5.030 2.460 5.260 3.405 ;
        RECT  5.010 0.635 5.240 1.410 ;
        RECT  4.660 3.175 5.030 3.405 ;
        RECT  4.660 0.635 5.010 0.865 ;
        RECT  4.800 1.760 4.975 2.100 ;
        RECT  4.570 1.760 4.800 2.735 ;
        RECT  4.295 2.495 4.570 2.735 ;
        RECT  4.065 2.495 4.295 3.220 ;
        RECT  2.825 2.990 4.065 3.220 ;
        RECT  3.195 0.520 3.445 2.755 ;
        RECT  1.845 0.520 3.195 0.760 ;
        RECT  3.105 2.525 3.195 2.755 ;
        RECT  2.585 1.000 2.825 3.220 ;
        RECT  2.345 1.000 2.585 1.240 ;
        RECT  2.345 2.670 2.585 2.910 ;
        RECT  2.075 1.680 2.315 2.360 ;
        RECT  1.845 2.130 2.075 2.775 ;
        RECT  1.625 0.520 1.845 1.415 ;
        RECT  0.470 2.545 1.845 2.775 ;
        RECT  1.605 0.520 1.625 1.980 ;
        RECT  1.385 1.175 1.605 1.980 ;
        RECT  0.380 0.560 0.480 0.900 ;
        RECT  0.380 2.545 0.470 3.440 ;
        RECT  0.140 0.560 0.380 3.440 ;
    END
END XOR3D1BWP7T

MACRO XOR3D2BWP7T
    CLASS CORE ;
    FOREIGN XOR3D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.080 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.125 0.970 9.380 3.075 ;
        RECT  9.100 0.490 9.125 3.385 ;
        RECT  8.895 0.490 9.100 1.305 ;
        RECT  8.895 2.795 9.100 3.385 ;
        END
    END Z
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 1.210 8.260 2.150 ;
        RECT  7.965 1.210 7.980 1.875 ;
        RECT  7.650 1.535 7.965 1.875 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4365 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.650 1.100 1.030 2.100 ;
        RECT  0.590 1.590 0.650 1.930 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 1.210 4.340 1.590 ;
        RECT  3.500 1.210 3.780 2.000 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 -0.235 10.080 0.235 ;
        RECT  9.615 -0.235 9.845 1.195 ;
        RECT  8.280 -0.235 9.615 0.235 ;
        RECT  7.940 -0.235 8.280 0.900 ;
        RECT  5.305 -0.235 7.940 0.235 ;
        RECT  5.075 -0.235 5.305 0.795 ;
        RECT  3.960 -0.235 5.075 0.235 ;
        RECT  3.580 -0.235 3.960 0.670 ;
        RECT  1.265 -0.235 3.580 0.235 ;
        RECT  0.885 -0.235 1.265 0.825 ;
        RECT  0.000 -0.235 0.885 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.845 3.685 10.080 4.155 ;
        RECT  9.615 2.255 9.845 4.155 ;
        RECT  8.345 3.685 9.615 4.155 ;
        RECT  7.885 3.250 8.345 4.155 ;
        RECT  5.390 3.685 7.885 4.155 ;
        RECT  5.050 3.225 5.390 4.155 ;
        RECT  4.130 3.685 5.050 4.155 ;
        RECT  3.790 3.340 4.130 4.155 ;
        RECT  1.290 3.685 3.790 4.155 ;
        RECT  0.910 3.250 1.290 4.155 ;
        RECT  0.000 3.685 0.910 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.720 1.735 8.870 1.975 ;
        RECT  8.490 1.735 8.720 2.610 ;
        RECT  8.290 2.380 8.490 2.610 ;
        RECT  8.060 2.380 8.290 3.020 ;
        RECT  6.885 2.790 8.060 3.020 ;
        RECT  7.350 2.330 7.560 2.560 ;
        RECT  7.350 1.020 7.520 1.250 ;
        RECT  7.115 0.465 7.350 2.560 ;
        RECT  5.840 0.465 7.115 0.695 ;
        RECT  6.655 0.950 6.885 3.020 ;
        RECT  6.380 0.950 6.655 1.180 ;
        RECT  6.500 2.300 6.655 2.530 ;
        RECT  5.850 3.225 6.470 3.455 ;
        RECT  6.195 1.410 6.425 1.970 ;
        RECT  5.960 1.740 6.195 1.970 ;
        RECT  5.730 1.740 5.960 2.410 ;
        RECT  5.620 2.765 5.850 3.455 ;
        RECT  5.610 0.465 5.840 1.255 ;
        RECT  4.840 2.180 5.730 2.410 ;
        RECT  4.700 2.765 5.620 2.995 ;
        RECT  5.500 1.025 5.610 1.255 ;
        RECT  5.260 1.025 5.500 1.950 ;
        RECT  4.610 0.560 4.840 2.535 ;
        RECT  4.360 2.765 4.700 3.315 ;
        RECT  4.300 0.560 4.610 0.790 ;
        RECT  4.290 2.295 4.610 2.535 ;
        RECT  2.765 2.765 4.360 2.995 ;
        RECT  3.230 2.305 3.360 2.535 ;
        RECT  2.995 0.875 3.230 2.535 ;
        RECT  2.920 0.875 2.995 1.105 ;
        RECT  2.690 0.465 2.920 1.105 ;
        RECT  1.750 3.225 2.820 3.455 ;
        RECT  2.535 1.335 2.765 2.995 ;
        RECT  1.725 0.465 2.690 0.695 ;
        RECT  2.460 1.335 2.535 1.565 ;
        RECT  2.260 2.525 2.535 2.755 ;
        RECT  2.120 0.925 2.460 1.565 ;
        RECT  1.965 1.800 2.305 2.140 ;
        RECT  1.735 1.800 1.965 2.560 ;
        RECT  1.520 2.790 1.750 3.455 ;
        RECT  0.360 2.330 1.735 2.560 ;
        RECT  1.495 0.465 1.725 1.385 ;
        RECT  0.625 2.790 1.520 3.020 ;
        RECT  1.265 1.155 1.495 1.770 ;
        RECT  0.395 2.790 0.625 3.370 ;
        RECT  0.360 0.540 0.480 0.880 ;
        RECT  0.130 0.540 0.360 2.560 ;
    END
END XOR3D2BWP7T

MACRO XOR4D0BWP7T
    CLASS CORE ;
    FOREIGN XOR4D0BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 0.5688 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 0.765 8.260 2.535 ;
        RECT  7.880 0.765 7.980 0.995 ;
        RECT  7.880 2.295 7.980 2.535 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.795 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.2133 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 1.600 9.205 1.960 ;
        RECT  8.540 1.210 8.820 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.210 12.180 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 -0.235 12.880 0.235 ;
        RECT  11.695 -0.235 11.930 0.980 ;
        RECT  9.040 -0.235 11.695 0.235 ;
        RECT  8.660 -0.235 9.040 0.970 ;
        RECT  5.495 -0.235 8.660 0.235 ;
        RECT  5.265 -0.235 5.495 1.225 ;
        RECT  4.130 -0.235 5.265 0.235 ;
        RECT  3.790 -0.235 4.130 0.915 ;
        RECT  1.185 -0.235 3.790 0.235 ;
        RECT  0.955 -0.235 1.185 0.980 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 3.685 12.880 4.155 ;
        RECT  11.695 3.025 11.930 4.155 ;
        RECT  8.980 3.685 11.695 4.155 ;
        RECT  8.615 3.445 8.980 4.155 ;
        RECT  5.495 3.685 8.615 4.155 ;
        RECT  5.265 2.710 5.495 4.155 ;
        RECT  4.130 3.685 5.265 4.155 ;
        RECT  3.790 3.455 4.130 4.155 ;
        RECT  1.185 3.685 3.790 4.155 ;
        RECT  0.955 2.980 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.410 0.670 12.650 3.230 ;
        RECT  11.500 2.510 12.410 2.750 ;
        RECT  11.270 2.035 11.500 2.750 ;
        RECT  11.235 0.465 11.465 1.755 ;
        RECT  10.690 2.035 11.270 2.275 ;
        RECT  9.770 0.465 11.235 0.695 ;
        RECT  10.460 1.820 10.690 2.275 ;
        RECT  10.230 0.945 10.505 1.185 ;
        RECT  10.230 2.585 10.505 2.815 ;
        RECT  10.000 0.945 10.230 2.995 ;
        RECT  7.445 2.765 10.000 2.995 ;
        RECT  9.540 0.465 9.770 2.530 ;
        RECT  9.400 0.725 9.540 0.955 ;
        RECT  9.405 2.300 9.540 2.530 ;
        RECT  6.915 3.225 7.860 3.455 ;
        RECT  7.375 0.545 7.510 0.805 ;
        RECT  7.375 2.510 7.445 2.995 ;
        RECT  7.145 0.545 7.375 2.995 ;
        RECT  5.965 0.545 7.145 0.785 ;
        RECT  6.685 1.015 6.915 3.455 ;
        RECT  6.400 1.015 6.685 1.255 ;
        RECT  6.440 2.550 6.685 2.780 ;
        RECT  6.225 1.555 6.455 2.285 ;
        RECT  4.925 2.055 6.225 2.285 ;
        RECT  5.730 0.545 5.965 1.685 ;
        RECT  5.725 0.545 5.730 1.825 ;
        RECT  5.495 1.455 5.725 1.825 ;
        RECT  4.695 1.020 4.925 2.995 ;
        RECT  4.490 1.020 4.695 1.250 ;
        RECT  4.490 2.765 4.695 2.995 ;
        RECT  4.290 1.720 4.465 2.060 ;
        RECT  4.060 1.720 4.290 2.640 ;
        RECT  3.995 2.400 4.060 2.640 ;
        RECT  3.755 2.400 3.995 3.225 ;
        RECT  2.800 2.985 3.755 3.225 ;
        RECT  3.260 2.525 3.405 2.755 ;
        RECT  3.260 0.680 3.390 0.910 ;
        RECT  3.030 0.465 3.260 2.755 ;
        RECT  1.645 0.465 3.030 0.695 ;
        RECT  2.570 0.945 2.800 3.225 ;
        RECT  2.290 0.945 2.570 1.180 ;
        RECT  2.345 2.470 2.570 2.810 ;
        RECT  2.105 1.800 2.340 2.140 ;
        RECT  1.875 1.800 2.105 2.670 ;
        RECT  0.465 2.430 1.875 2.670 ;
        RECT  1.415 0.465 1.645 1.950 ;
        RECT  1.330 1.610 1.415 1.950 ;
        RECT  0.235 0.640 0.465 3.250 ;
    END
END XOR4D0BWP7T

MACRO XOR4D1BWP7T
    CLASS CORE ;
    FOREIGN XOR4D1BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.880 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.0312 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.980 0.765 8.260 2.535 ;
        RECT  7.880 0.765 7.980 0.995 ;
        RECT  7.880 2.295 7.980 2.535 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.795 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 1.600 9.205 1.960 ;
        RECT  8.540 1.210 8.820 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.900 1.210 12.180 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 -0.235 12.880 0.235 ;
        RECT  11.695 -0.235 11.930 0.980 ;
        RECT  9.040 -0.235 11.695 0.235 ;
        RECT  8.660 -0.235 9.040 0.970 ;
        RECT  5.495 -0.235 8.660 0.235 ;
        RECT  5.265 -0.235 5.495 1.225 ;
        RECT  4.130 -0.235 5.265 0.235 ;
        RECT  3.790 -0.235 4.130 0.915 ;
        RECT  1.185 -0.235 3.790 0.235 ;
        RECT  0.955 -0.235 1.185 0.980 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.930 3.685 12.880 4.155 ;
        RECT  11.695 3.025 11.930 4.155 ;
        RECT  8.980 3.685 11.695 4.155 ;
        RECT  8.615 3.445 8.980 4.155 ;
        RECT  5.495 3.685 8.615 4.155 ;
        RECT  5.265 2.710 5.495 4.155 ;
        RECT  4.130 3.685 5.265 4.155 ;
        RECT  3.790 3.455 4.130 4.155 ;
        RECT  1.185 3.685 3.790 4.155 ;
        RECT  0.955 2.980 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.410 0.670 12.650 3.230 ;
        RECT  11.500 2.510 12.410 2.750 ;
        RECT  11.270 2.035 11.500 2.750 ;
        RECT  11.235 0.465 11.465 1.755 ;
        RECT  10.690 2.035 11.270 2.275 ;
        RECT  9.770 0.465 11.235 0.695 ;
        RECT  10.460 1.820 10.690 2.275 ;
        RECT  10.230 0.945 10.505 1.185 ;
        RECT  10.230 2.585 10.505 2.815 ;
        RECT  10.000 0.945 10.230 2.995 ;
        RECT  7.445 2.765 10.000 2.995 ;
        RECT  9.540 0.465 9.770 2.530 ;
        RECT  9.400 0.725 9.540 0.955 ;
        RECT  9.405 2.300 9.540 2.530 ;
        RECT  6.915 3.225 7.860 3.455 ;
        RECT  7.375 0.545 7.510 0.805 ;
        RECT  7.375 2.510 7.445 2.995 ;
        RECT  7.145 0.545 7.375 2.995 ;
        RECT  5.965 0.545 7.145 0.785 ;
        RECT  6.685 1.015 6.915 3.455 ;
        RECT  6.400 1.015 6.685 1.255 ;
        RECT  6.440 2.550 6.685 2.780 ;
        RECT  6.225 1.555 6.455 2.285 ;
        RECT  4.925 2.055 6.225 2.285 ;
        RECT  5.730 0.545 5.965 1.685 ;
        RECT  5.725 0.545 5.730 1.825 ;
        RECT  5.495 1.455 5.725 1.825 ;
        RECT  4.695 1.020 4.925 2.995 ;
        RECT  4.490 1.020 4.695 1.250 ;
        RECT  4.490 2.765 4.695 2.995 ;
        RECT  4.290 1.720 4.465 2.060 ;
        RECT  4.060 1.720 4.290 2.640 ;
        RECT  3.995 2.400 4.060 2.640 ;
        RECT  3.755 2.400 3.995 3.225 ;
        RECT  2.800 2.985 3.755 3.225 ;
        RECT  3.260 2.525 3.405 2.755 ;
        RECT  3.260 0.680 3.390 0.910 ;
        RECT  3.030 0.465 3.260 2.755 ;
        RECT  1.645 0.465 3.030 0.695 ;
        RECT  2.570 0.945 2.800 3.225 ;
        RECT  2.290 0.945 2.570 1.180 ;
        RECT  2.345 2.470 2.570 2.810 ;
        RECT  2.105 1.800 2.340 2.140 ;
        RECT  1.875 1.800 2.105 2.670 ;
        RECT  0.465 2.430 1.875 2.670 ;
        RECT  1.415 0.465 1.645 1.950 ;
        RECT  1.330 1.610 1.415 1.950 ;
        RECT  0.235 0.640 0.465 3.250 ;
    END
END XOR4D1BWP7T

MACRO XOR4D2BWP7T
    CLASS CORE ;
    FOREIGN XOR4D2BWP7T 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.440 BY 3.920 ;
    SYMMETRY x y ;
    SITE core7T ;
    PIN Z
        ANTENNADIFFAREA 1.2798 ;
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.820 0.765 8.940 0.995 ;
        RECT  8.820 2.325 8.940 2.560 ;
        RECT  8.540 0.765 8.820 2.560 ;
        END
    END Z
    PIN A4
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.210 0.980 2.150 ;
        END
    END A4
    PIN A3
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.500 1.210 3.795 2.150 ;
        END
    END A3
    PIN A2
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.655 1.210 9.940 2.150 ;
        END
    END A2
    PIN A1
        ANTENNAGATEAREA 0.4266 ;
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.460 1.210 12.740 2.150 ;
        END
    END A1
    PIN VSS
        DIRECTION INOUT ;
        USE ground ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.490 -0.235 13.440 0.235 ;
        RECT  12.255 -0.235 12.490 0.980 ;
        RECT  9.700 -0.235 12.255 0.235 ;
        RECT  9.320 -0.235 9.700 0.970 ;
        RECT  8.220 -0.235 9.320 0.235 ;
        RECT  7.880 -0.235 8.220 0.725 ;
        RECT  5.495 -0.235 7.880 0.235 ;
        RECT  5.265 -0.235 5.495 1.225 ;
        RECT  4.130 -0.235 5.265 0.235 ;
        RECT  3.790 -0.235 4.130 0.915 ;
        RECT  1.185 -0.235 3.790 0.235 ;
        RECT  0.955 -0.235 1.185 0.980 ;
        RECT  0.000 -0.235 0.955 0.235 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE power ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.490 3.685 13.440 4.155 ;
        RECT  12.255 3.025 12.490 4.155 ;
        RECT  9.700 3.685 12.255 4.155 ;
        RECT  9.335 3.250 9.700 4.155 ;
        RECT  8.220 3.685 9.335 4.155 ;
        RECT  7.880 3.250 8.220 4.155 ;
        RECT  5.495 3.685 7.880 4.155 ;
        RECT  5.265 2.710 5.495 4.155 ;
        RECT  4.130 3.685 5.265 4.155 ;
        RECT  3.790 3.455 4.130 4.155 ;
        RECT  1.185 3.685 3.790 4.155 ;
        RECT  0.955 2.980 1.185 4.155 ;
        RECT  0.000 3.685 0.955 4.155 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.970 0.670 13.210 3.230 ;
        RECT  12.060 2.510 12.970 2.750 ;
        RECT  11.830 2.035 12.060 2.750 ;
        RECT  12.025 1.195 12.055 1.755 ;
        RECT  11.825 0.465 12.025 1.755 ;
        RECT  11.385 2.035 11.830 2.275 ;
        RECT  11.795 0.465 11.825 1.425 ;
        RECT  10.465 0.465 11.795 0.695 ;
        RECT  11.155 1.820 11.385 2.275 ;
        RECT  10.925 0.945 11.200 1.185 ;
        RECT  10.925 2.585 11.200 2.815 ;
        RECT  10.695 0.945 10.925 3.020 ;
        RECT  8.140 2.790 10.695 3.020 ;
        RECT  10.235 0.465 10.465 2.560 ;
        RECT  10.095 0.725 10.235 0.955 ;
        RECT  10.100 2.330 10.235 2.560 ;
        RECT  7.900 1.090 8.140 3.020 ;
        RECT  7.470 1.090 7.900 1.330 ;
        RECT  7.235 2.465 7.900 2.805 ;
        RECT  6.915 1.600 7.655 1.940 ;
        RECT  7.230 0.545 7.470 1.330 ;
        RECT  5.965 0.545 7.230 0.785 ;
        RECT  6.685 1.015 6.915 2.780 ;
        RECT  6.400 1.015 6.685 1.255 ;
        RECT  6.440 2.550 6.685 2.780 ;
        RECT  6.225 1.555 6.455 2.285 ;
        RECT  4.925 2.055 6.225 2.285 ;
        RECT  5.730 0.545 5.965 1.685 ;
        RECT  5.725 0.545 5.730 1.825 ;
        RECT  5.495 1.455 5.725 1.825 ;
        RECT  4.695 1.020 4.925 2.995 ;
        RECT  4.490 1.020 4.695 1.250 ;
        RECT  4.490 2.765 4.695 2.995 ;
        RECT  4.290 1.720 4.465 2.060 ;
        RECT  4.060 1.720 4.290 2.640 ;
        RECT  3.995 2.400 4.060 2.640 ;
        RECT  3.755 2.400 3.995 3.225 ;
        RECT  2.800 2.985 3.755 3.225 ;
        RECT  3.260 2.525 3.405 2.755 ;
        RECT  3.260 0.680 3.390 0.910 ;
        RECT  3.030 0.465 3.260 2.755 ;
        RECT  1.645 0.465 3.030 0.695 ;
        RECT  2.570 0.945 2.800 3.225 ;
        RECT  2.290 0.945 2.570 1.180 ;
        RECT  2.345 2.470 2.570 2.810 ;
        RECT  2.105 1.800 2.340 2.140 ;
        RECT  1.875 1.800 2.105 2.670 ;
        RECT  0.465 2.430 1.875 2.670 ;
        RECT  1.415 0.465 1.645 1.950 ;
        RECT  1.330 1.610 1.415 1.950 ;
        RECT  0.235 0.640 0.465 3.250 ;
    END
END XOR4D2BWP7T

END LIBRARY
